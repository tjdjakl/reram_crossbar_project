magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< pwell >>
rect 467 350 491 401
<< metal1 >>
rect 0 911 876 918
rect 0 859 52 911
rect 104 859 116 911
rect 168 859 180 911
rect 232 859 244 911
rect 296 859 308 911
rect 360 859 516 911
rect 568 859 580 911
rect 632 859 644 911
rect 696 859 708 911
rect 760 859 772 911
rect 824 859 876 911
rect 0 852 876 859
rect 0 842 66 852
rect 0 790 7 842
rect 59 790 66 842
rect 0 778 66 790
rect 0 726 7 778
rect 59 726 66 778
rect 0 714 66 726
rect 0 662 7 714
rect 59 662 66 714
rect 0 650 66 662
rect 0 598 7 650
rect 59 598 66 650
rect 0 586 66 598
rect 0 534 7 586
rect 59 534 66 586
rect 0 384 66 534
rect 0 332 7 384
rect 59 332 66 384
rect 0 320 66 332
rect 0 268 7 320
rect 59 268 66 320
rect 0 256 66 268
rect 0 204 7 256
rect 59 204 66 256
rect 0 192 66 204
rect 0 140 7 192
rect 59 140 66 192
rect 0 128 66 140
rect 0 76 7 128
rect 59 76 66 128
rect 113 491 141 824
rect 169 519 197 852
rect 225 491 253 824
rect 281 519 309 852
rect 337 491 365 824
rect 411 818 465 824
rect 411 766 412 818
rect 464 766 465 818
rect 411 754 465 766
rect 411 702 412 754
rect 464 702 465 754
rect 411 690 465 702
rect 411 638 412 690
rect 464 638 465 690
rect 411 626 465 638
rect 411 574 412 626
rect 464 574 465 626
rect 411 562 465 574
rect 411 510 412 562
rect 464 510 465 562
rect 411 491 465 510
rect 511 491 539 824
rect 567 519 595 852
rect 623 491 651 824
rect 679 519 707 852
rect 810 842 876 852
rect 735 491 763 824
rect 113 485 763 491
rect 113 433 119 485
rect 171 433 183 485
rect 235 433 247 485
rect 299 433 311 485
rect 363 433 513 485
rect 565 433 577 485
rect 629 433 641 485
rect 693 433 705 485
rect 757 433 763 485
rect 113 427 763 433
rect 113 94 141 427
rect 0 66 66 76
rect 169 66 197 399
rect 225 94 253 427
rect 281 66 309 399
rect 337 94 365 427
rect 411 408 465 427
rect 411 356 412 408
rect 464 356 465 408
rect 411 344 465 356
rect 411 292 412 344
rect 464 292 465 344
rect 411 280 465 292
rect 411 228 412 280
rect 464 228 465 280
rect 411 216 465 228
rect 411 164 412 216
rect 464 164 465 216
rect 411 152 465 164
rect 411 100 412 152
rect 464 100 465 152
rect 411 94 465 100
rect 511 94 539 427
rect 567 66 595 399
rect 623 94 651 427
rect 679 66 707 399
rect 735 94 763 427
rect 810 790 817 842
rect 869 790 876 842
rect 810 778 876 790
rect 810 726 817 778
rect 869 726 876 778
rect 810 714 876 726
rect 810 662 817 714
rect 869 662 876 714
rect 810 650 876 662
rect 810 598 817 650
rect 869 598 876 650
rect 810 586 876 598
rect 810 534 817 586
rect 869 534 876 586
rect 810 384 876 534
rect 810 332 817 384
rect 869 332 876 384
rect 810 320 876 332
rect 810 268 817 320
rect 869 268 876 320
rect 810 256 876 268
rect 810 204 817 256
rect 869 204 876 256
rect 810 192 876 204
rect 810 140 817 192
rect 869 140 876 192
rect 810 128 876 140
rect 810 76 817 128
rect 869 76 876 128
rect 810 66 876 76
rect 0 59 876 66
rect 0 7 52 59
rect 104 7 116 59
rect 168 7 180 59
rect 232 7 244 59
rect 296 7 308 59
rect 360 7 516 59
rect 568 7 580 59
rect 632 7 644 59
rect 696 7 708 59
rect 760 7 772 59
rect 824 7 876 59
rect 0 0 876 7
<< via1 >>
rect 52 859 104 911
rect 116 859 168 911
rect 180 859 232 911
rect 244 859 296 911
rect 308 859 360 911
rect 516 859 568 911
rect 580 859 632 911
rect 644 859 696 911
rect 708 859 760 911
rect 772 859 824 911
rect 7 790 59 842
rect 7 726 59 778
rect 7 662 59 714
rect 7 598 59 650
rect 7 534 59 586
rect 7 332 59 384
rect 7 268 59 320
rect 7 204 59 256
rect 7 140 59 192
rect 7 76 59 128
rect 412 766 464 818
rect 412 702 464 754
rect 412 638 464 690
rect 412 574 464 626
rect 412 510 464 562
rect 119 433 171 485
rect 183 433 235 485
rect 247 433 299 485
rect 311 433 363 485
rect 513 433 565 485
rect 577 433 629 485
rect 641 433 693 485
rect 705 433 757 485
rect 412 356 464 408
rect 412 292 464 344
rect 412 228 464 280
rect 412 164 464 216
rect 412 100 464 152
rect 817 790 869 842
rect 817 726 869 778
rect 817 662 869 714
rect 817 598 869 650
rect 817 534 869 586
rect 817 332 869 384
rect 817 268 869 320
rect 817 204 869 256
rect 817 140 869 192
rect 817 76 869 128
rect 52 7 104 59
rect 116 7 168 59
rect 180 7 232 59
rect 244 7 296 59
rect 308 7 360 59
rect 516 7 568 59
rect 580 7 632 59
rect 644 7 696 59
rect 708 7 760 59
rect 772 7 824 59
<< metal2 >>
rect 0 911 383 918
rect 0 859 52 911
rect 104 859 116 911
rect 168 859 180 911
rect 232 859 244 911
rect 296 859 308 911
rect 360 859 383 911
rect 0 852 383 859
rect 0 842 66 852
rect 0 790 7 842
rect 59 790 66 842
rect 411 824 465 918
rect 493 911 876 918
rect 493 859 516 911
rect 568 859 580 911
rect 632 859 644 911
rect 696 859 708 911
rect 760 859 772 911
rect 824 859 876 911
rect 493 852 876 859
rect 810 842 876 852
rect 94 818 782 824
rect 94 796 412 818
rect 0 778 66 790
rect 0 726 7 778
rect 59 768 66 778
rect 59 740 383 768
rect 411 766 412 796
rect 464 796 782 818
rect 464 766 465 796
rect 810 790 817 842
rect 869 790 876 842
rect 810 778 876 790
rect 810 768 817 778
rect 411 754 465 766
rect 59 726 66 740
rect 0 714 66 726
rect 0 662 7 714
rect 59 662 66 714
rect 411 712 412 754
rect 94 702 412 712
rect 464 712 465 754
rect 493 740 817 768
rect 810 726 817 740
rect 869 726 876 778
rect 810 714 876 726
rect 464 702 782 712
rect 94 690 782 702
rect 94 684 412 690
rect 0 656 66 662
rect 0 650 383 656
rect 0 598 7 650
rect 59 628 383 650
rect 411 638 412 684
rect 464 684 782 690
rect 464 638 465 684
rect 810 662 817 714
rect 869 662 876 714
rect 810 656 876 662
rect 59 598 66 628
rect 411 626 465 638
rect 493 650 876 656
rect 493 628 817 650
rect 411 600 412 626
rect 0 586 66 598
rect 0 534 7 586
rect 59 544 66 586
rect 94 574 412 600
rect 464 600 465 626
rect 464 574 782 600
rect 94 572 782 574
rect 810 598 817 628
rect 869 598 876 650
rect 810 586 876 598
rect 411 562 465 572
rect 59 534 383 544
rect 0 516 383 534
rect 411 510 412 562
rect 464 510 465 562
rect 810 544 817 586
rect 493 534 817 544
rect 869 534 876 586
rect 493 516 876 534
rect 411 488 465 510
rect 0 485 876 488
rect 0 433 119 485
rect 171 433 183 485
rect 235 433 247 485
rect 299 433 311 485
rect 363 433 513 485
rect 565 433 577 485
rect 629 433 641 485
rect 693 433 705 485
rect 757 433 876 485
rect 0 430 876 433
rect 411 408 465 430
rect 0 384 383 402
rect 0 332 7 384
rect 59 374 383 384
rect 59 332 66 374
rect 411 356 412 408
rect 464 356 465 408
rect 493 384 876 402
rect 493 374 817 384
rect 411 346 465 356
rect 0 320 66 332
rect 0 268 7 320
rect 59 290 66 320
rect 94 344 782 346
rect 94 318 412 344
rect 411 292 412 318
rect 464 318 782 344
rect 810 332 817 374
rect 869 332 876 384
rect 810 320 876 332
rect 464 292 465 318
rect 59 268 383 290
rect 0 262 383 268
rect 411 280 465 292
rect 810 290 817 320
rect 0 256 66 262
rect 0 204 7 256
rect 59 204 66 256
rect 411 234 412 280
rect 94 228 412 234
rect 464 234 465 280
rect 493 268 817 290
rect 869 268 876 320
rect 493 262 876 268
rect 810 256 876 262
rect 464 228 782 234
rect 94 216 782 228
rect 94 206 412 216
rect 0 192 66 204
rect 0 140 7 192
rect 59 178 66 192
rect 59 150 383 178
rect 411 164 412 206
rect 464 206 782 216
rect 464 164 465 206
rect 810 204 817 256
rect 869 204 876 256
rect 810 192 876 204
rect 810 178 817 192
rect 411 152 465 164
rect 59 140 66 150
rect 0 128 66 140
rect 0 76 7 128
rect 59 76 66 128
rect 411 122 412 152
rect 94 100 412 122
rect 464 122 465 152
rect 493 150 817 178
rect 810 140 817 150
rect 869 140 876 192
rect 810 128 876 140
rect 464 100 782 122
rect 94 94 782 100
rect 0 66 66 76
rect 0 59 383 66
rect 0 7 52 59
rect 104 7 116 59
rect 168 7 180 59
rect 232 7 244 59
rect 296 7 308 59
rect 360 7 383 59
rect 0 0 383 7
rect 411 0 465 94
rect 810 76 817 128
rect 869 76 876 128
rect 810 66 876 76
rect 493 59 876 66
rect 493 7 516 59
rect 568 7 580 59
rect 632 7 644 59
rect 696 7 708 59
rect 760 7 772 59
rect 824 7 876 59
rect 493 0 876 7
<< labels >>
flabel metal2 s 291 634 317 649 0 FreeSans 400 0 0 0 C0
port 2 nsew
flabel metal2 s 420 755 458 792 0 FreeSans 400 0 0 0 C1
port 3 nsew
flabel pwell s 467 350 491 401 0 FreeSans 200 0 0 0 SUB
port 4 nsew
<< properties >>
string GDS_END 169568
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 160160
<< end >>
