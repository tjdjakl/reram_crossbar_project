magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 978 203
rect 30 -17 64 21
<< locali >>
rect 17 199 66 323
rect 638 323 704 425
rect 806 323 872 425
rect 638 289 872 323
rect 638 170 714 289
rect 748 204 995 255
rect 638 127 995 170
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 391 69 493
rect 103 425 175 527
rect 17 357 175 391
rect 100 265 175 357
rect 215 345 257 493
rect 291 379 357 527
rect 391 345 425 493
rect 459 379 531 527
rect 565 459 995 493
rect 565 345 599 459
rect 215 311 599 345
rect 738 357 772 459
rect 906 289 995 459
rect 100 199 604 265
rect 100 165 139 199
rect 17 131 139 165
rect 207 131 604 165
rect 17 51 69 131
rect 103 17 169 97
rect 207 51 241 131
rect 275 17 341 97
rect 375 51 409 131
rect 443 17 511 97
rect 547 93 604 131
rect 547 51 995 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 748 204 995 255 6 A
port 1 nsew signal input
rlabel locali s 17 199 66 323 6 TE
port 2 nsew signal input
rlabel metal1 s 0 -48 1012 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 978 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1050 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 638 127 995 170 6 Z
port 7 nsew signal output
rlabel locali s 638 170 714 289 6 Z
port 7 nsew signal output
rlabel locali s 638 289 872 323 6 Z
port 7 nsew signal output
rlabel locali s 806 323 872 425 6 Z
port 7 nsew signal output
rlabel locali s 638 323 704 425 6 Z
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1012 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2038900
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2030936
<< end >>
