magic
tech sky130B
magscale 1 2
timestamp 1700618825
<< metal1 >>
rect 5058 4914 5258 4944
rect 5058 4774 5082 4914
rect 5246 4774 5258 4914
rect 10846 4804 10856 4944
rect 11020 4804 11030 4944
rect 14492 4860 14502 5000
rect 14666 4860 14676 5000
rect 5058 4744 5258 4774
rect 6904 1444 7098 2578
rect 4014 1232 4214 1270
rect 6904 1244 7192 1444
rect 4014 1072 4024 1232
rect 4174 1072 4214 1232
rect 9770 1110 9780 1268
rect 9938 1110 9948 1268
rect 4014 1070 4214 1072
rect 12682 992 12872 2558
rect 16330 2552 16530 2752
rect 13420 1150 13620 1350
rect 5388 736 5588 936
rect 6096 756 6296 956
rect 12680 852 12690 992
rect 12854 852 12872 992
rect 12682 842 12872 852
<< via1 >>
rect 5082 4774 5246 4914
rect 10856 4804 11020 4944
rect 14502 4860 14666 5000
rect 4024 1072 4174 1232
rect 9780 1110 9938 1268
rect 12690 852 12854 992
<< metal2 >>
rect 14502 5000 14666 5010
rect 5092 4944 14502 4994
rect 5092 4924 10856 4944
rect 5082 4914 10856 4924
rect 5246 4804 10856 4914
rect 11020 4860 14502 4944
rect 11020 4850 14666 4860
rect 11020 4804 14610 4850
rect 5246 4774 14610 4804
rect 5082 4766 14610 4774
rect 5082 4764 5246 4766
rect 9780 1268 9938 1278
rect 4024 1232 4174 1242
rect 9780 1100 9938 1110
rect 4024 1062 4174 1072
rect 12690 992 12854 1002
rect 11190 926 11340 936
rect 5400 910 5568 920
rect 12854 854 14964 988
rect 12690 842 12854 852
rect 11190 770 11340 780
rect 5400 724 5568 734
<< via2 >>
rect 4024 1072 4174 1232
rect 9780 1110 9938 1268
rect 5400 734 5568 910
rect 11190 780 11340 926
<< metal3 >>
rect 9770 1268 9948 1273
rect 4014 1232 4184 1237
rect 9770 1232 9780 1268
rect 4014 1072 4024 1232
rect 4174 1110 9780 1232
rect 9938 1110 9948 1268
rect 4174 1105 9948 1110
rect 4174 1072 9922 1105
rect 4014 1067 9922 1072
rect 4058 1050 9922 1067
rect 11180 926 11350 931
rect 5390 910 5578 915
rect 11180 910 11190 926
rect 5390 734 5400 910
rect 5568 780 11190 910
rect 11340 780 11350 926
rect 5568 775 11350 780
rect 5568 734 11344 775
rect 5390 729 5578 734
use invOpAmp  invOpAmp_0
timestamp 1700618825
transform 1 0 8592 0 1 260
box -1422 340 4296 9042
use TIA_04  TIA_04_1
timestamp 1700618825
transform 1 0 3512 0 1 164
box 240 340 3596 9210
use oneBitADC  x4
timestamp 1700618825
transform 1 0 12234 0 1 312
box 656 288 4296 4810
<< labels >>
flabel metal1 4014 1070 4214 1270 0 FreeSans 256 0 0 0 VSSneg
port 3 nsew
flabel metal1 5388 736 5588 936 0 FreeSans 256 0 0 0 Gnd
port 4 nsew
flabel metal1 13420 1150 13620 1350 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 16330 2552 16530 2752 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 5058 4744 5258 4944 0 FreeSans 256 0 0 0 VDD18
port 1 nsew
flabel metal1 6096 756 6296 956 0 FreeSans 256 0 0 0 Vin
port 0 nsew
<< end >>
