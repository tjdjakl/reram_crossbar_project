magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 42 201 1525 203
rect 42 23 1831 201
rect 42 21 339 23
rect 836 21 1028 23
rect 1440 21 1831 23
rect 42 17 63 21
rect 29 -17 63 17
<< locali >>
rect 164 409 214 493
rect 109 288 214 409
rect 109 185 172 288
rect 109 132 210 185
rect 160 70 210 132
rect 464 199 591 265
rect 1429 289 1545 323
rect 1429 199 1463 289
rect 1593 215 1675 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 60 443 130 527
rect 248 443 315 527
rect 352 447 671 481
rect 714 447 795 481
rect 829 447 895 527
rect 962 455 1581 489
rect 1663 455 1730 527
rect 352 409 386 447
rect 761 413 795 447
rect 962 413 996 455
rect 248 375 386 409
rect 466 379 727 413
rect 761 379 996 413
rect 248 265 282 375
rect 329 307 659 341
rect 242 199 282 265
rect 248 173 282 199
rect 248 139 362 173
rect 60 17 126 93
rect 244 17 294 105
rect 328 85 362 139
rect 396 119 430 307
rect 625 265 659 307
rect 693 339 727 379
rect 693 305 799 339
rect 742 275 799 305
rect 625 199 680 265
rect 486 131 708 165
rect 570 85 640 91
rect 328 51 640 85
rect 674 85 708 131
rect 742 119 776 275
rect 833 241 867 379
rect 913 289 996 343
rect 810 207 867 241
rect 810 85 844 207
rect 674 51 844 85
rect 878 17 912 173
rect 948 83 996 289
rect 1031 119 1065 421
rect 1099 178 1133 455
rect 1764 421 1823 493
rect 1171 323 1254 409
rect 1361 387 1823 421
rect 1171 289 1327 323
rect 1174 199 1259 254
rect 1099 165 1143 178
rect 1099 144 1182 165
rect 1109 131 1182 144
rect 1031 97 1075 119
rect 1031 53 1114 97
rect 1148 64 1182 131
rect 1216 126 1259 199
rect 1293 85 1327 289
rect 1361 119 1395 387
rect 1726 375 1823 387
rect 1579 299 1743 341
rect 1709 265 1743 299
rect 1497 189 1559 255
rect 1709 199 1755 265
rect 1497 146 1538 189
rect 1709 181 1743 199
rect 1595 150 1743 181
rect 1587 147 1743 150
rect 1429 85 1522 93
rect 1293 51 1522 85
rect 1587 59 1645 147
rect 1789 117 1823 375
rect 1679 17 1713 113
rect 1763 51 1823 117
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< obsm1 >>
rect 753 320 811 329
rect 1213 320 1271 329
rect 753 292 1271 320
rect 753 283 811 292
rect 1213 283 1271 292
rect 937 184 995 193
rect 1213 184 1271 193
rect 1489 184 1547 193
rect 937 156 1547 184
rect 937 147 995 156
rect 1213 147 1271 156
rect 1489 147 1547 156
rect 1029 116 1087 125
rect 1581 116 1639 125
rect 1029 88 1639 116
rect 1029 79 1087 88
rect 1581 79 1639 88
<< labels >>
rlabel locali s 1593 215 1675 265 6 A
port 1 nsew signal input
rlabel locali s 1429 199 1463 289 6 B
port 2 nsew signal input
rlabel locali s 1429 289 1545 323 6 B
port 2 nsew signal input
rlabel locali s 464 199 591 265 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 1840 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 42 17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1440 21 1831 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 836 21 1028 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 42 21 339 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 42 23 1831 201 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 42 201 1525 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1878 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1840 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 160 70 210 132 6 X
port 8 nsew signal output
rlabel locali s 109 132 210 185 6 X
port 8 nsew signal output
rlabel locali s 109 185 172 288 6 X
port 8 nsew signal output
rlabel locali s 109 288 214 409 6 X
port 8 nsew signal output
rlabel locali s 164 409 214 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1840 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 685594
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 673288
<< end >>
