magic
tech sky130B
magscale 1 2
timestamp 1700618825
<< locali >>
rect 990 1578 1692 1638
rect 990 1438 1224 1578
rect 1680 1438 1692 1578
rect 990 1286 1692 1438
rect 990 584 1146 1286
rect 1534 584 1692 1286
rect 990 580 1112 584
rect 1568 580 1692 584
rect 990 382 1108 384
rect 1568 382 1690 384
rect 990 -186 1146 382
rect 1534 -186 1690 382
rect 990 -244 1690 -186
rect 990 -384 1224 -244
rect 1680 -384 1690 -244
rect 990 -444 1690 -384
<< viali >>
rect 1224 1438 1680 1578
rect 1224 -384 1680 -244
<< metal1 >>
rect 990 1578 1692 1638
rect 990 1438 1224 1578
rect 1680 1438 1692 1578
rect 990 1300 1692 1438
rect 1204 950 1262 1300
rect 1318 780 1358 1178
rect 1438 1004 1462 1006
rect 896 502 1096 576
rect 1314 502 1360 780
rect 896 432 1360 502
rect 896 376 1096 432
rect 1314 192 1360 432
rect 1412 502 1462 1004
rect 1580 502 1780 572
rect 1412 432 1780 502
rect 1204 -154 1262 118
rect 1320 -48 1354 192
rect 1412 70 1462 432
rect 1580 372 1780 432
rect 990 -244 1690 -154
rect 990 -384 1224 -244
rect 1680 -384 1690 -244
rect 990 -444 1690 -384
use sky130_fd_pr__nfet_g5v0d10v5_6XHARQ  XM1 ~/Project/magic
timestamp 1700618825
transform 1 0 1338 0 1 99
box -278 -333 278 333
use sky130_fd_pr__pfet_g5v0d10v5_7EBZY6  XM2 ~/Project/magic
timestamp 1700618825
transform 1 0 1338 0 1 949
box -308 -447 308 447
<< labels >>
flabel metal1 1002 1414 1202 1614 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 1000 -420 1200 -220 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 896 376 1096 576 0 FreeSans 256 0 0 0 Vin
port 0 nsew
flabel metal1 1580 372 1780 572 0 FreeSans 256 0 0 0 Vout
port 3 nsew
<< end >>
