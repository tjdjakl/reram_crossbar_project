magic
tech sky130B
magscale 1 2
timestamp 1700618825
<< locali >>
rect 468 2058 2898 2070
rect 468 1918 526 2058
rect 1274 2054 2898 2058
rect 1274 1918 1508 2054
rect 2854 1918 2898 2054
rect 468 456 638 1918
rect 736 1758 2898 1918
rect 736 456 1410 1758
rect 468 136 1410 456
rect 222 -1540 348 -28
rect 1000 -428 1136 -28
rect 1294 -174 1410 136
rect 2748 -174 2898 1758
rect 1000 -530 1410 -428
rect 1000 -694 1058 -530
rect 1000 -892 1150 -694
rect 1244 -892 1410 -530
rect 1000 -1348 1410 -892
rect 1000 -1540 1138 -1348
rect 222 -1564 1138 -1540
rect 1288 -1540 1410 -1348
rect 2748 -1540 2868 -428
rect 1288 -1564 2868 -1540
rect 222 -1702 2868 -1564
rect 222 -1808 442 -1702
rect 2820 -1808 2868 -1702
rect 222 -1832 2868 -1808
<< viali >>
rect 526 1918 1274 2058
rect 1508 1918 2854 2054
rect 638 456 736 1918
rect 1058 -694 1244 -530
rect 1150 -892 1244 -694
rect 1138 -1564 1288 -1348
rect 442 -1808 2820 -1702
<< metal1 >>
rect 468 2058 2898 2070
rect 468 1918 526 2058
rect 1274 2054 2898 2058
rect 1274 1918 1508 2054
rect 2854 1918 2898 2054
rect 468 1758 638 1918
rect 586 1462 638 1758
rect 736 1758 2898 1918
rect 736 1462 774 1758
rect 576 1178 586 1462
rect 774 1178 784 1462
rect 586 456 638 1178
rect 736 456 774 1178
rect 586 -164 774 456
rect 1348 24 1520 218
rect 402 -1352 412 -994
rect 474 -1352 484 -994
rect 612 -1474 756 -164
rect 1348 -242 1442 24
rect 1660 2 1812 1690
rect 1926 1164 1936 1476
rect 1996 1164 2006 1476
rect 2038 26 2210 220
rect 1654 -22 1834 2
rect 1654 -38 1664 -22
rect 1628 -148 1664 -38
rect 1834 -148 1844 -22
rect 1628 -242 1834 -148
rect 1348 -348 1834 -242
rect 2038 -254 2132 26
rect 2342 2 2508 1690
rect 2610 1162 2620 1474
rect 2680 1162 2690 1474
rect 2324 -20 2528 2
rect 2324 -146 2344 -20
rect 2514 -146 2528 -20
rect 2324 -196 2528 -146
rect 3138 -254 3338 -222
rect 886 -522 1216 -520
rect 886 -530 1280 -522
rect 886 -694 1058 -530
rect 886 -706 1150 -694
rect 1130 -892 1150 -706
rect 1244 -892 1280 -530
rect 1348 -688 1442 -348
rect 2038 -380 3338 -254
rect 1348 -866 1524 -688
rect 1130 -996 1280 -892
rect 1114 -1332 1292 -996
rect 1102 -1348 1322 -1332
rect 1102 -1540 1138 -1348
rect 228 -1564 1138 -1540
rect 1288 -1540 1322 -1348
rect 1658 -1428 1824 -530
rect 2038 -686 2132 -380
rect 3138 -422 3338 -380
rect 2038 -864 2214 -686
rect 1924 -1350 1934 -992
rect 1996 -1350 2006 -992
rect 2348 -1428 2514 -530
rect 2612 -1346 2622 -988
rect 2684 -1346 2694 -988
rect 1628 -1500 1638 -1428
rect 1850 -1500 1860 -1428
rect 2328 -1500 2338 -1428
rect 2550 -1500 2560 -1428
rect 1288 -1564 2862 -1540
rect 228 -1702 2862 -1564
rect 228 -1808 442 -1702
rect 2820 -1808 2862 -1702
rect 228 -1824 2862 -1808
rect 1610 -1954 1852 -1922
rect 1610 -2158 1646 -1954
rect 1840 -2158 1852 -1954
rect 2324 -1932 2566 -1910
rect 2324 -2136 2338 -1932
rect 2532 -2136 2566 -1932
rect 2324 -2146 2566 -2136
<< via1 >>
rect 586 1178 638 1462
rect 638 1178 736 1462
rect 736 1178 774 1462
rect 412 -1352 474 -994
rect 1936 1164 1996 1476
rect 1664 -148 1834 -22
rect 2620 1162 2680 1474
rect 2344 -146 2514 -20
rect 1934 -1350 1996 -992
rect 2622 -1346 2684 -988
rect 1638 -1500 1850 -1428
rect 2338 -1500 2550 -1428
rect 1646 -2158 1840 -1954
rect 2338 -2136 2532 -1932
<< metal2 >>
rect 1936 1476 1996 1486
rect 586 1462 774 1472
rect 774 1178 1936 1462
rect 586 1168 774 1178
rect 2620 1474 2680 1484
rect 1996 1178 2620 1462
rect 1936 1154 1996 1164
rect 2620 1152 2680 1162
rect 1664 -20 1834 -12
rect 2344 -20 2514 -10
rect 1664 -22 2344 -20
rect 1834 -146 2344 -22
rect 2514 -146 2530 -20
rect 1834 -148 2530 -146
rect 1664 -158 1834 -148
rect 2344 -156 2514 -148
rect 412 -994 474 -984
rect 1934 -992 1996 -982
rect 474 -1332 1934 -1004
rect 412 -1362 474 -1352
rect 2622 -988 2684 -978
rect 1996 -1332 2622 -1004
rect 1934 -1360 1996 -1350
rect 2622 -1356 2684 -1346
rect 1638 -1428 1850 -1418
rect 1638 -1510 1850 -1500
rect 2338 -1428 2550 -1418
rect 2338 -1510 2550 -1500
rect 1656 -1944 1826 -1510
rect 2352 -1922 2512 -1510
rect 2338 -1932 2532 -1922
rect 1646 -1954 1840 -1944
rect 2338 -2146 2532 -2136
rect 1646 -2168 1840 -2158
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XM5 ~/Project/magic
timestamp 1700618825
transform 1 0 1736 0 1 809
box -396 -1019 396 1019
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XM6
timestamp 1700618825
transform 1 0 2422 0 1 809
box -396 -1019 396 1019
use sky130_fd_pr__nfet_01v8_AHRV9L  XM16 ~/Project/magic
timestamp 1700618825
transform 1 0 2422 0 1 -1002
box -396 -610 396 610
use sky130_fd_pr__nfet_01v8_lvt_XVWV9B  XM17 ~/Project/magic
timestamp 1700618825
transform 1 0 674 0 1 -802
box -396 -810 396 810
use sky130_fd_pr__nfet_01v8_AHRV9L  XM23
timestamp 1700618825
transform 1 0 1736 0 1 -1002
box -396 -610 396 610
<< labels >>
flabel metal1 3138 -422 3338 -222 0 FreeSans 256 0 0 0 Vout
port 5 nsew
flabel metal1 228 -1824 428 -1624 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 2334 -2122 2534 -1922 0 FreeSans 256 0 0 0 Vminus
port 4 nsew
flabel metal1 1630 -2142 1830 -1942 0 FreeSans 256 0 0 0 Vplus
port 3 nsew
flabel metal1 1294 1868 1494 2068 0 FreeSans 256 0 0 0 VCC
port 1 nsew
<< end >>
