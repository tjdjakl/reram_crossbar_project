magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 98 157 1318 203
rect 1 21 1318 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 176 47 206 177
rect 370 47 400 177
rect 454 47 484 177
rect 538 47 568 177
rect 622 47 652 177
rect 706 47 736 177
rect 790 47 820 177
rect 874 47 904 177
rect 958 47 988 177
rect 1042 47 1072 177
rect 1126 47 1156 177
rect 1210 47 1240 177
<< scpmoshvt >>
rect 79 297 109 425
rect 176 297 206 497
rect 370 297 400 497
rect 454 297 484 497
rect 538 297 568 497
rect 622 297 652 497
rect 706 297 736 497
rect 790 297 820 497
rect 874 297 904 497
rect 958 297 988 497
rect 1042 297 1072 497
rect 1126 297 1156 497
rect 1210 297 1240 497
<< ndiff >>
rect 124 131 176 177
rect 27 111 79 131
rect 27 77 35 111
rect 69 77 79 111
rect 27 47 79 77
rect 109 97 176 131
rect 109 63 119 97
rect 153 63 176 97
rect 109 47 176 63
rect 206 165 258 177
rect 206 131 216 165
rect 250 131 258 165
rect 206 97 258 131
rect 206 63 216 97
rect 250 63 258 97
rect 206 47 258 63
rect 318 165 370 177
rect 318 131 326 165
rect 360 131 370 165
rect 318 97 370 131
rect 318 63 326 97
rect 360 63 370 97
rect 318 47 370 63
rect 400 97 454 177
rect 400 63 410 97
rect 444 63 454 97
rect 400 47 454 63
rect 484 165 538 177
rect 484 131 494 165
rect 528 131 538 165
rect 484 97 538 131
rect 484 63 494 97
rect 528 63 538 97
rect 484 47 538 63
rect 568 97 622 177
rect 568 63 578 97
rect 612 63 622 97
rect 568 47 622 63
rect 652 165 706 177
rect 652 131 662 165
rect 696 131 706 165
rect 652 97 706 131
rect 652 63 662 97
rect 696 63 706 97
rect 652 47 706 63
rect 736 97 790 177
rect 736 63 746 97
rect 780 63 790 97
rect 736 47 790 63
rect 820 165 874 177
rect 820 131 830 165
rect 864 131 874 165
rect 820 97 874 131
rect 820 63 830 97
rect 864 63 874 97
rect 820 47 874 63
rect 904 97 958 177
rect 904 63 914 97
rect 948 63 958 97
rect 904 47 958 63
rect 988 165 1042 177
rect 988 131 998 165
rect 1032 131 1042 165
rect 988 97 1042 131
rect 988 63 998 97
rect 1032 63 1042 97
rect 988 47 1042 63
rect 1072 97 1126 177
rect 1072 63 1082 97
rect 1116 63 1126 97
rect 1072 47 1126 63
rect 1156 165 1210 177
rect 1156 131 1166 165
rect 1200 131 1210 165
rect 1156 97 1210 131
rect 1156 63 1166 97
rect 1200 63 1210 97
rect 1156 47 1210 63
rect 1240 97 1292 177
rect 1240 63 1250 97
rect 1284 63 1292 97
rect 1240 47 1292 63
<< pdiff >>
rect 124 425 176 497
rect 27 411 79 425
rect 27 377 35 411
rect 69 377 79 411
rect 27 343 79 377
rect 27 309 35 343
rect 69 309 79 343
rect 27 297 79 309
rect 109 407 176 425
rect 109 373 119 407
rect 153 373 176 407
rect 109 297 176 373
rect 206 479 258 497
rect 206 445 216 479
rect 250 445 258 479
rect 206 411 258 445
rect 206 377 216 411
rect 250 377 258 411
rect 206 343 258 377
rect 206 309 216 343
rect 250 309 258 343
rect 206 297 258 309
rect 318 479 370 497
rect 318 445 326 479
rect 360 445 370 479
rect 318 411 370 445
rect 318 377 326 411
rect 360 377 370 411
rect 318 343 370 377
rect 318 309 326 343
rect 360 309 370 343
rect 318 297 370 309
rect 400 485 454 497
rect 400 451 410 485
rect 444 451 454 485
rect 400 417 454 451
rect 400 383 410 417
rect 444 383 454 417
rect 400 297 454 383
rect 484 479 538 497
rect 484 445 494 479
rect 528 445 538 479
rect 484 411 538 445
rect 484 377 494 411
rect 528 377 538 411
rect 484 343 538 377
rect 484 309 494 343
rect 528 309 538 343
rect 484 297 538 309
rect 568 485 622 497
rect 568 451 578 485
rect 612 451 622 485
rect 568 417 622 451
rect 568 383 578 417
rect 612 383 622 417
rect 568 297 622 383
rect 652 479 706 497
rect 652 445 662 479
rect 696 445 706 479
rect 652 411 706 445
rect 652 377 662 411
rect 696 377 706 411
rect 652 343 706 377
rect 652 309 662 343
rect 696 309 706 343
rect 652 297 706 309
rect 736 485 790 497
rect 736 451 746 485
rect 780 451 790 485
rect 736 417 790 451
rect 736 383 746 417
rect 780 383 790 417
rect 736 297 790 383
rect 820 479 874 497
rect 820 445 830 479
rect 864 445 874 479
rect 820 411 874 445
rect 820 377 830 411
rect 864 377 874 411
rect 820 343 874 377
rect 820 309 830 343
rect 864 309 874 343
rect 820 297 874 309
rect 904 485 958 497
rect 904 451 914 485
rect 948 451 958 485
rect 904 417 958 451
rect 904 383 914 417
rect 948 383 958 417
rect 904 297 958 383
rect 988 479 1042 497
rect 988 445 998 479
rect 1032 445 1042 479
rect 988 411 1042 445
rect 988 377 998 411
rect 1032 377 1042 411
rect 988 343 1042 377
rect 988 309 998 343
rect 1032 309 1042 343
rect 988 297 1042 309
rect 1072 485 1126 497
rect 1072 451 1082 485
rect 1116 451 1126 485
rect 1072 417 1126 451
rect 1072 383 1082 417
rect 1116 383 1126 417
rect 1072 297 1126 383
rect 1156 479 1210 497
rect 1156 445 1166 479
rect 1200 445 1210 479
rect 1156 411 1210 445
rect 1156 377 1166 411
rect 1200 377 1210 411
rect 1156 343 1210 377
rect 1156 309 1166 343
rect 1200 309 1210 343
rect 1156 297 1210 309
rect 1240 485 1292 497
rect 1240 451 1250 485
rect 1284 451 1292 485
rect 1240 417 1292 451
rect 1240 383 1250 417
rect 1284 383 1292 417
rect 1240 297 1292 383
<< ndiffc >>
rect 35 77 69 111
rect 119 63 153 97
rect 216 131 250 165
rect 216 63 250 97
rect 326 131 360 165
rect 326 63 360 97
rect 410 63 444 97
rect 494 131 528 165
rect 494 63 528 97
rect 578 63 612 97
rect 662 131 696 165
rect 662 63 696 97
rect 746 63 780 97
rect 830 131 864 165
rect 830 63 864 97
rect 914 63 948 97
rect 998 131 1032 165
rect 998 63 1032 97
rect 1082 63 1116 97
rect 1166 131 1200 165
rect 1166 63 1200 97
rect 1250 63 1284 97
<< pdiffc >>
rect 35 377 69 411
rect 35 309 69 343
rect 119 373 153 407
rect 216 445 250 479
rect 216 377 250 411
rect 216 309 250 343
rect 326 445 360 479
rect 326 377 360 411
rect 326 309 360 343
rect 410 451 444 485
rect 410 383 444 417
rect 494 445 528 479
rect 494 377 528 411
rect 494 309 528 343
rect 578 451 612 485
rect 578 383 612 417
rect 662 445 696 479
rect 662 377 696 411
rect 662 309 696 343
rect 746 451 780 485
rect 746 383 780 417
rect 830 445 864 479
rect 830 377 864 411
rect 830 309 864 343
rect 914 451 948 485
rect 914 383 948 417
rect 998 445 1032 479
rect 998 377 1032 411
rect 998 309 1032 343
rect 1082 451 1116 485
rect 1082 383 1116 417
rect 1166 445 1200 479
rect 1166 377 1200 411
rect 1166 309 1200 343
rect 1250 451 1284 485
rect 1250 383 1284 417
<< poly >>
rect 176 497 206 523
rect 370 497 400 523
rect 454 497 484 523
rect 538 497 568 523
rect 622 497 652 523
rect 706 497 736 523
rect 790 497 820 523
rect 874 497 904 523
rect 958 497 988 523
rect 1042 497 1072 523
rect 1126 497 1156 523
rect 1210 497 1240 523
rect 79 425 109 451
rect 79 265 109 297
rect 176 265 206 297
rect 22 249 109 265
rect 22 215 38 249
rect 72 215 109 249
rect 22 199 109 215
rect 161 249 218 265
rect 161 215 174 249
rect 208 215 218 249
rect 161 199 218 215
rect 370 259 400 297
rect 454 259 484 297
rect 538 259 568 297
rect 370 249 568 259
rect 370 215 410 249
rect 444 215 478 249
rect 512 215 568 249
rect 370 205 568 215
rect 79 131 109 199
rect 176 177 206 199
rect 370 177 400 205
rect 454 177 484 205
rect 538 177 568 205
rect 622 259 652 297
rect 706 259 736 297
rect 790 259 820 297
rect 874 259 904 297
rect 958 259 988 297
rect 1042 259 1072 297
rect 1126 259 1156 297
rect 1210 259 1240 297
rect 622 249 1240 259
rect 622 215 646 249
rect 680 215 714 249
rect 748 215 782 249
rect 816 215 850 249
rect 884 215 918 249
rect 952 215 986 249
rect 1020 215 1240 249
rect 622 205 1240 215
rect 622 177 652 205
rect 706 177 736 205
rect 790 177 820 205
rect 874 177 904 205
rect 958 177 988 205
rect 1042 177 1072 205
rect 1126 177 1156 205
rect 1210 177 1240 205
rect 79 21 109 47
rect 176 21 206 47
rect 370 21 400 47
rect 454 21 484 47
rect 538 21 568 47
rect 622 21 652 47
rect 706 21 736 47
rect 790 21 820 47
rect 874 21 904 47
rect 958 21 988 47
rect 1042 21 1072 47
rect 1126 21 1156 47
rect 1210 21 1240 47
<< polycont >>
rect 38 215 72 249
rect 174 215 208 249
rect 410 215 444 249
rect 478 215 512 249
rect 646 215 680 249
rect 714 215 748 249
rect 782 215 816 249
rect 850 215 884 249
rect 918 215 952 249
rect 986 215 1020 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 19 411 85 432
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 119 407 153 527
rect 119 357 153 373
rect 200 479 276 493
rect 200 445 216 479
rect 250 445 276 479
rect 200 411 276 445
rect 200 377 216 411
rect 250 377 276 411
rect 19 309 35 343
rect 69 323 85 343
rect 200 343 276 377
rect 69 309 156 323
rect 200 309 216 343
rect 250 309 276 343
rect 19 289 156 309
rect 122 265 156 289
rect 22 249 88 255
rect 22 215 38 249
rect 72 215 88 249
rect 122 249 208 265
rect 122 215 174 249
rect 122 199 208 215
rect 242 255 276 309
rect 310 479 376 493
rect 310 445 326 479
rect 360 445 376 479
rect 310 411 376 445
rect 310 377 326 411
rect 360 377 376 411
rect 310 343 376 377
rect 410 485 444 527
rect 410 417 444 451
rect 410 357 444 383
rect 478 479 544 493
rect 478 445 494 479
rect 528 445 544 479
rect 478 411 544 445
rect 478 377 494 411
rect 528 377 544 411
rect 310 309 326 343
rect 360 323 376 343
rect 478 343 544 377
rect 578 485 612 527
rect 578 417 612 451
rect 578 357 612 383
rect 646 479 712 493
rect 646 445 662 479
rect 696 445 712 479
rect 646 411 712 445
rect 646 377 662 411
rect 696 377 712 411
rect 478 323 494 343
rect 360 309 494 323
rect 528 323 544 343
rect 646 343 712 377
rect 746 485 780 527
rect 746 417 780 451
rect 746 367 780 383
rect 814 479 880 493
rect 814 445 830 479
rect 864 445 880 479
rect 814 411 880 445
rect 814 377 830 411
rect 864 377 880 411
rect 528 309 612 323
rect 310 289 612 309
rect 646 309 662 343
rect 696 323 712 343
rect 814 343 880 377
rect 914 485 948 527
rect 914 417 948 451
rect 914 367 948 383
rect 982 479 1048 493
rect 982 445 998 479
rect 1032 445 1048 479
rect 982 411 1048 445
rect 982 377 998 411
rect 1032 377 1048 411
rect 814 323 830 343
rect 696 309 830 323
rect 864 323 880 343
rect 982 343 1048 377
rect 1082 485 1116 527
rect 1082 417 1116 451
rect 1082 367 1116 383
rect 1150 479 1216 493
rect 1150 445 1166 479
rect 1200 445 1216 479
rect 1150 411 1216 445
rect 1150 377 1166 411
rect 1200 377 1216 411
rect 982 323 998 343
rect 864 309 998 323
rect 1032 323 1048 343
rect 1150 343 1216 377
rect 1250 485 1284 527
rect 1250 417 1284 451
rect 1250 367 1284 383
rect 1150 323 1166 343
rect 1032 309 1166 323
rect 1200 323 1216 343
rect 1200 309 1363 323
rect 646 289 1363 309
rect 578 255 612 289
rect 242 249 544 255
rect 242 215 410 249
rect 444 215 478 249
rect 512 215 544 249
rect 578 249 1072 255
rect 578 215 646 249
rect 680 215 714 249
rect 748 215 782 249
rect 816 215 850 249
rect 884 215 918 249
rect 952 215 986 249
rect 1020 215 1072 249
rect 122 181 156 199
rect 19 147 156 181
rect 242 165 276 215
rect 578 181 612 215
rect 1287 181 1363 289
rect 19 111 85 147
rect 200 131 216 165
rect 250 131 276 165
rect 19 77 35 111
rect 69 77 85 111
rect 19 52 85 77
rect 119 97 153 113
rect 119 17 153 63
rect 200 97 276 131
rect 200 63 216 97
rect 250 63 276 97
rect 200 52 276 63
rect 310 165 612 181
rect 310 131 326 165
rect 360 147 494 165
rect 360 131 376 147
rect 310 97 376 131
rect 478 131 494 147
rect 528 147 612 165
rect 646 165 1363 181
rect 528 131 544 147
rect 310 63 326 97
rect 360 63 376 97
rect 310 52 376 63
rect 410 97 444 113
rect 410 17 444 63
rect 478 97 544 131
rect 646 131 662 165
rect 696 147 830 165
rect 696 131 712 147
rect 478 63 494 97
rect 528 63 544 97
rect 478 52 544 63
rect 578 97 612 113
rect 578 17 612 63
rect 646 97 712 131
rect 814 131 830 147
rect 864 147 998 165
rect 864 131 880 147
rect 646 63 662 97
rect 696 63 712 97
rect 646 52 712 63
rect 746 97 780 113
rect 746 17 780 63
rect 814 97 880 131
rect 982 131 998 147
rect 1032 147 1166 165
rect 1032 131 1048 147
rect 814 63 830 97
rect 864 63 880 97
rect 814 52 880 63
rect 914 97 948 113
rect 914 17 948 63
rect 982 97 1048 131
rect 1150 131 1166 147
rect 1200 147 1363 165
rect 1200 131 1216 147
rect 982 63 998 97
rect 1032 63 1048 97
rect 982 52 1048 63
rect 1082 97 1116 113
rect 1082 17 1116 63
rect 1150 97 1216 131
rect 1150 63 1166 97
rect 1200 63 1216 97
rect 1150 52 1216 63
rect 1250 97 1284 113
rect 1250 17 1284 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1317 221 1351 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 1317 289 1351 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 bufbuf_8
rlabel metal1 s 0 -48 1380 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1380 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_END 3258950
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3248478
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 34.500 0.000 
<< end >>
