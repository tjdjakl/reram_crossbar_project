magic
tech sky130B
magscale 1 2
timestamp 1700618825
<< pwell >>
rect -253 -710 253 710
<< psubdiff >>
rect -217 640 -121 674
rect 121 640 217 674
rect -217 578 -183 640
rect 183 578 217 640
rect -217 -640 -183 -578
rect 183 -640 217 -578
rect -217 -674 -121 -640
rect 121 -674 217 -640
<< psubdiffcont >>
rect -121 640 121 674
rect -217 -578 -183 578
rect 183 -578 217 578
rect -121 -674 121 -640
<< poly >>
rect -87 -494 -21 -114
rect -87 -528 -71 -494
rect -37 -528 -21 -494
rect -87 -544 -21 -528
rect 21 -494 87 -114
rect 21 -528 37 -494
rect 71 -528 87 -494
rect 21 -544 87 -528
<< polycont >>
rect -71 -528 -37 -494
rect 37 -528 71 -494
<< npolyres >>
rect -87 478 87 544
rect -87 -114 -21 478
rect 21 -114 87 478
<< locali >>
rect -217 640 -121 674
rect 121 640 217 674
rect -217 578 -183 640
rect 183 578 217 640
rect -87 -528 -71 -494
rect -37 -528 -21 -494
rect 21 -528 37 -494
rect 71 -528 87 -494
rect -217 -640 -183 -578
rect 183 -640 217 -578
rect -217 -674 -121 -640
rect 121 -674 217 -640
<< properties >>
string FIXED_BBOX -200 -657 200 657
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.33 l 2.77 m 1 nx 2 wmin 0.330 lmin 1.650 rho 48.2 val 915.8 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 1 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
