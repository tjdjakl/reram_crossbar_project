magic
tech sky130B
magscale 1 2
timestamp 1700618825
<< pwell >>
rect -253 -1053 253 1053
<< psubdiff >>
rect -217 983 -121 1017
rect 121 983 217 1017
rect -217 921 -183 983
rect 183 921 217 983
rect -217 -983 -183 -921
rect 183 -983 217 -921
rect -217 -1017 -121 -983
rect 121 -1017 217 -983
<< psubdiffcont >>
rect -121 983 121 1017
rect -217 -921 -183 921
rect 183 -921 217 921
rect -121 -1017 121 -983
<< poly >>
rect -87 -837 -21 -457
rect -87 -871 -71 -837
rect -37 -871 -21 -837
rect -87 -887 -21 -871
rect 21 -837 87 -457
rect 21 -871 37 -837
rect 71 -871 87 -837
rect 21 -887 87 -871
<< polycont >>
rect -71 -871 -37 -837
rect 37 -871 71 -837
<< npolyres >>
rect -87 821 87 887
rect -87 -457 -21 821
rect 21 -457 87 821
<< locali >>
rect -217 983 -121 1017
rect 121 983 217 1017
rect -217 921 -183 983
rect 183 921 217 983
rect -87 -871 -71 -837
rect -37 -871 -21 -837
rect 21 -871 37 -837
rect 71 -871 87 -837
rect -217 -983 -183 -921
rect 183 -983 217 -921
rect -217 -1017 -121 -983
rect 121 -1017 217 -983
<< properties >>
string FIXED_BBOX -200 -1000 200 1000
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w .33 l 6.2 m 1 nx 2 wmin 0.330 lmin 1.650 rho 48.2 val 1.917k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 1 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
