magic
tech sky130B
magscale 1 2
timestamp 1700640585
<< locali >>
rect -842 2714 90 2716
rect -140 2403 90 2714
rect -185 2376 94 2403
rect -140 1656 90 2376
rect 804 1684 1034 2716
rect -142 900 88 1460
rect -142 820 100 900
rect -142 632 88 820
rect -842 600 88 632
rect 806 600 1026 1432
<< metal1 >>
rect -842 2714 94 2716
rect -830 2490 -630 2690
rect -140 2403 94 2714
rect 800 2406 1056 2716
rect -924 2244 -724 2298
rect -924 2142 -894 2244
rect -772 2142 -724 2244
rect 32 2210 42 2284
rect 134 2210 144 2284
rect 946 2192 956 2272
rect 1074 2192 1084 2272
rect -924 2098 -724 2142
rect -936 1594 -736 1652
rect -936 1494 -900 1594
rect -764 1494 -736 1594
rect 1624 1590 1824 1644
rect -936 1452 -736 1494
rect -232 1492 -222 1590
rect -94 1492 -84 1590
rect 14 1506 24 1568
rect 142 1506 152 1568
rect 702 1474 712 1576
rect 852 1474 862 1576
rect 964 1490 974 1572
rect 1104 1490 1114 1572
rect 1624 1488 1654 1590
rect 1794 1488 1824 1590
rect 1624 1444 1824 1488
rect -924 1134 -724 1186
rect -924 1032 -890 1134
rect -768 1032 -724 1134
rect -924 986 -724 1032
rect 28 996 38 1076
rect 156 996 166 1076
rect 954 1024 964 1096
rect 1056 1024 1066 1096
rect -832 656 -632 856
rect -142 820 -140 882
rect -142 632 88 820
rect -842 600 88 632
rect 806 600 1038 882
<< via1 >>
rect -894 2142 -772 2244
rect 42 2210 134 2284
rect 956 2192 1074 2272
rect -900 1494 -764 1594
rect -222 1492 -94 1590
rect 24 1506 142 1568
rect 712 1474 852 1576
rect 974 1490 1104 1572
rect 1654 1488 1794 1590
rect -890 1032 -768 1134
rect 38 996 156 1076
rect 964 1024 1056 1096
<< metal2 >>
rect 42 2284 134 2294
rect -894 2244 -772 2254
rect -894 2132 -772 2142
rect -222 2210 42 2284
rect -900 1594 -764 1604
rect -900 1484 -764 1494
rect -222 1590 -94 2210
rect 42 2200 134 2210
rect 956 2272 1074 2282
rect 956 2182 1074 2192
rect 712 1806 1738 1930
rect 24 1568 142 1578
rect 24 1496 142 1506
rect 712 1576 852 1806
rect 1646 1596 1738 1806
rect 1646 1590 1794 1596
rect -222 1384 -94 1492
rect 974 1572 1104 1582
rect 1646 1546 1654 1590
rect 974 1480 1104 1490
rect 1654 1478 1794 1488
rect 712 1464 852 1474
rect -222 1260 1056 1384
rect -890 1134 -768 1144
rect 964 1096 1056 1260
rect -890 1022 -768 1032
rect 38 1076 156 1086
rect 964 1014 1056 1024
rect 38 986 156 996
<< via2 >>
rect -894 2142 -772 2244
rect -900 1494 -764 1594
rect 956 2192 1074 2272
rect 24 1506 142 1568
rect 974 1490 1104 1572
rect -890 1032 -768 1134
rect 38 996 156 1076
<< metal3 >>
rect 946 2272 1084 2277
rect -904 2244 -762 2249
rect -904 2142 -894 2244
rect -772 2142 -22 2244
rect 946 2192 956 2272
rect 1074 2192 1084 2272
rect 946 2187 1084 2192
rect -904 2137 -762 2142
rect -142 1798 -22 2142
rect -142 1710 104 1798
rect -910 1594 -754 1599
rect -910 1494 -900 1594
rect -764 1494 -754 1594
rect 26 1573 104 1710
rect 14 1568 152 1573
rect 14 1506 24 1568
rect 142 1506 152 1568
rect 14 1501 152 1506
rect 964 1572 1114 1577
rect -910 1489 -754 1494
rect 964 1490 974 1572
rect 1104 1490 1114 1572
rect 964 1485 1114 1490
rect 1004 1422 1098 1485
rect -890 1324 1098 1422
rect -890 1139 -768 1324
rect -900 1134 -758 1139
rect -900 1032 -890 1134
rect -768 1032 -758 1134
rect -900 1027 -758 1032
rect 28 1076 166 1081
rect 28 996 38 1076
rect 156 996 166 1076
rect 28 991 166 996
<< via3 >>
rect 956 2192 1074 2272
rect -900 1494 -764 1594
rect 38 996 156 1076
<< metal4 >>
rect 955 2272 1075 2273
rect 955 2192 956 2272
rect 1074 2192 1075 2272
rect 955 2191 1075 2192
rect -901 1594 -763 1595
rect -901 1494 -900 1594
rect -764 1592 -763 1594
rect 960 1592 1036 2191
rect -764 1494 1036 1592
rect -901 1493 -763 1494
rect 36 1077 154 1494
rect 36 1076 157 1077
rect 36 1026 38 1076
rect 37 996 38 1026
rect 156 996 157 1076
rect 37 995 157 996
use TransmissionGate  x1
timestamp 1700624956
transform 1 0 -126 0 1 180
box 126 420 1016 2536
use TransmissionGate  x2
timestamp 1700624956
transform 1 0 808 0 1 180
box 126 420 1016 2536
use Inverter  x3
timestamp 1700618825
transform 1 0 -1832 0 1 1076
box 896 -444 1780 1638
<< labels >>
flabel metal1 -924 2098 -724 2298 0 FreeSans 256 0 0 0 A
port 0 nsew
flabel metal1 -924 986 -724 1186 0 FreeSans 256 0 0 0 B
port 1 nsew
flabel metal1 -936 1452 -736 1652 0 FreeSans 256 0 0 0 S
port 2 nsew
flabel metal1 -830 2490 -630 2690 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 -832 656 -632 856 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 1624 1444 1824 1644 0 FreeSans 256 0 0 0 OUT
port 5 nsew
<< end >>
