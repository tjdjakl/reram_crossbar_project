magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< poly >>
rect 264 10020 424 10036
rect 264 9986 293 10020
rect 327 9986 361 10020
rect 395 9986 424 10020
rect 264 9652 293 9686
rect 327 9652 361 9686
rect 395 9652 424 9686
rect 264 9636 424 9652
rect 520 10000 680 10016
rect 520 9966 549 10000
rect 583 9966 617 10000
rect 651 9966 680 10000
rect 520 9632 549 9666
rect 583 9632 617 9666
rect 651 9632 680 9666
rect 520 9616 680 9632
rect 264 9435 424 9451
rect 264 9401 293 9435
rect 327 9401 361 9435
rect 395 9401 424 9435
rect 264 9067 293 9101
rect 327 9067 361 9101
rect 395 9067 424 9101
rect 264 9051 424 9067
rect 520 9415 680 9431
rect 520 9381 549 9415
rect 583 9381 617 9415
rect 651 9381 680 9415
rect 520 9047 549 9081
rect 583 9047 617 9081
rect 651 9047 680 9081
rect 520 9031 680 9047
<< polycont >>
rect 293 9986 327 10020
rect 361 9986 395 10020
rect 293 9652 327 9686
rect 361 9652 395 9686
rect 549 9966 583 10000
rect 617 9966 651 10000
rect 549 9632 583 9666
rect 617 9632 651 9666
rect 293 9401 327 9435
rect 361 9401 395 9435
rect 293 9067 327 9101
rect 361 9067 395 9101
rect 549 9381 583 9415
rect 617 9381 651 9415
rect 549 9047 583 9081
rect 617 9047 651 9081
<< npolyres >>
rect 264 9686 424 9986
rect 520 9666 680 9966
rect 264 9101 424 9401
rect 520 9081 680 9381
<< locali >>
rect 277 9993 291 10099
rect 397 9993 411 10099
rect 277 9986 293 9993
rect 327 9986 361 9993
rect 395 9986 411 9993
rect 533 9994 547 10100
rect 653 9994 667 10100
rect 533 9966 549 9994
rect 583 9966 617 9994
rect 651 9966 667 9994
rect 277 9665 293 9686
rect 277 9631 291 9665
rect 327 9652 361 9686
rect 395 9665 411 9686
rect 325 9631 363 9652
rect 397 9631 411 9665
rect 277 9537 411 9631
rect 277 9431 291 9537
rect 397 9431 411 9537
rect 277 9401 293 9431
rect 327 9401 361 9431
rect 395 9401 411 9431
rect 533 9632 547 9666
rect 583 9632 617 9666
rect 653 9632 667 9666
rect 533 9548 667 9632
rect 533 9442 547 9548
rect 653 9442 667 9548
rect 533 9415 667 9442
rect 533 9381 549 9415
rect 583 9381 617 9415
rect 651 9381 667 9415
rect 277 9067 291 9101
rect 327 9067 361 9101
rect 397 9067 411 9101
rect 533 9047 547 9081
rect 583 9047 617 9081
rect 653 9047 667 9081
rect 327 8908 365 8942
rect 578 8772 616 8806
rect 325 7674 363 7708
rect 325 7566 363 7600
rect 325 6332 363 6366
rect 276 5434 410 6080
rect 276 5328 468 5434
<< viali >>
rect 291 10020 397 10099
rect 291 9993 293 10020
rect 293 9993 327 10020
rect 327 9993 361 10020
rect 361 9993 395 10020
rect 395 9993 397 10020
rect 547 10000 653 10100
rect 547 9994 549 10000
rect 549 9994 583 10000
rect 583 9994 617 10000
rect 617 9994 651 10000
rect 651 9994 653 10000
rect 291 9652 293 9665
rect 293 9652 325 9665
rect 363 9652 395 9665
rect 395 9652 397 9665
rect 291 9631 325 9652
rect 363 9631 397 9652
rect 291 9435 397 9537
rect 291 9431 293 9435
rect 293 9431 327 9435
rect 327 9431 361 9435
rect 361 9431 395 9435
rect 395 9431 397 9435
rect 547 9632 549 9666
rect 549 9632 581 9666
rect 619 9632 651 9666
rect 651 9632 653 9666
rect 547 9442 653 9548
rect 291 9067 293 9101
rect 293 9067 325 9101
rect 363 9067 395 9101
rect 395 9067 397 9101
rect 547 9047 549 9081
rect 549 9047 581 9081
rect 619 9047 651 9081
rect 651 9047 653 9081
rect 293 8908 327 8942
rect 365 8908 399 8942
rect 544 8772 578 8806
rect 616 8772 650 8806
rect 291 7674 325 7708
rect 363 7674 397 7708
rect 291 7566 325 7600
rect 363 7566 397 7600
rect 291 6332 325 6366
rect 363 6332 397 6366
rect 468 5328 646 5434
<< metal1 >>
tri 282 10218 342 10278 se
rect 342 10218 607 10278
tri 607 10218 667 10278 sw
tri 277 10213 282 10218 se
rect 282 10213 667 10218
rect 277 10150 667 10213
rect 277 10099 409 10150
tri 409 10123 436 10150 nw
tri 507 10123 534 10150 ne
rect 534 10123 667 10150
tri 534 10122 535 10123 ne
rect 277 9993 291 10099
rect 397 9993 409 10099
rect 277 9980 409 9993
rect 278 9978 408 9979
rect 277 9678 409 9978
rect 278 9677 408 9678
rect 277 9665 409 9676
rect 277 9631 291 9665
rect 325 9631 363 9665
rect 397 9631 409 9665
rect 277 9537 409 9631
rect 277 9431 291 9537
rect 397 9431 409 9537
rect 277 9420 409 9431
rect 278 9418 408 9419
rect 277 9118 409 9418
rect 278 9117 408 9118
rect 277 9101 409 9116
rect 277 9067 291 9101
rect 325 9067 363 9101
rect 397 9067 409 9101
rect 277 9064 409 9067
rect 535 10100 667 10123
rect 535 9994 547 10100
rect 653 9994 667 10100
rect 535 9980 667 9994
rect 536 9978 666 9979
rect 535 9678 667 9978
rect 536 9677 666 9678
rect 535 9666 667 9676
rect 535 9632 547 9666
rect 581 9632 619 9666
rect 653 9632 667 9666
rect 535 9548 667 9632
rect 535 9442 547 9548
rect 653 9442 667 9548
rect 535 9399 667 9442
rect 536 9397 666 9398
rect 535 9097 667 9397
rect 536 9096 666 9097
rect 535 9081 667 9095
tri 277 9062 279 9064 ne
rect 279 9062 409 9064
tri 409 9062 411 9064 sw
rect 279 8942 411 9062
rect 535 9047 547 9081
rect 581 9047 619 9081
rect 653 9047 667 9081
rect 535 9041 667 9047
rect 279 8908 293 8942
rect 327 8908 365 8942
rect 399 8908 411 8942
rect 279 8591 411 8908
rect 280 8589 410 8590
rect 279 8289 411 8589
rect 280 8288 410 8289
rect 279 7708 411 8287
rect 279 7674 291 7708
rect 325 7674 363 7708
rect 397 7674 411 7708
rect 279 7600 411 7674
rect 279 7566 291 7600
rect 325 7566 363 7600
rect 397 7566 411 7600
rect 279 7375 411 7566
rect 280 7373 410 7374
rect 532 8806 662 8812
rect 532 8772 544 8806
rect 578 8772 616 8806
rect 650 8772 662 8806
rect 280 7072 410 7073
rect 279 6860 411 7071
tri 411 6860 436 6885 sw
tri 507 6860 532 6885 se
rect 532 6860 662 8772
rect 279 6779 662 6860
rect 279 6366 409 6779
tri 409 6752 436 6779 nw
rect 279 6332 291 6366
rect 325 6332 363 6366
rect 397 6332 409 6366
rect 279 6326 409 6332
rect 456 5434 658 5440
rect 456 5328 468 5434
rect 646 5328 658 5434
rect 456 5322 658 5328
<< rmetal1 >>
rect 277 9979 409 9980
rect 277 9978 278 9979
rect 408 9978 409 9979
rect 277 9677 278 9678
rect 408 9677 409 9678
rect 277 9676 409 9677
rect 277 9419 409 9420
rect 277 9418 278 9419
rect 408 9418 409 9419
rect 277 9117 278 9118
rect 408 9117 409 9118
rect 277 9116 409 9117
rect 535 9979 667 9980
rect 535 9978 536 9979
rect 666 9978 667 9979
rect 535 9677 536 9678
rect 666 9677 667 9678
rect 535 9676 667 9677
rect 535 9398 667 9399
rect 535 9397 536 9398
rect 666 9397 667 9398
rect 535 9096 536 9097
rect 666 9096 667 9097
rect 535 9095 667 9096
rect 279 8590 411 8591
rect 279 8589 280 8590
rect 410 8589 411 8590
rect 279 8288 280 8289
rect 410 8288 411 8289
rect 279 8287 411 8288
rect 279 7374 411 7375
rect 279 7373 280 7374
rect 410 7373 411 7374
rect 279 7072 280 7073
rect 410 7072 411 7073
rect 279 7071 411 7072
use sky130_fd_io__gpio_ovtv2_res_weak_bentbigres  sky130_fd_io__gpio_ovtv2_res_weak_bentbigres_0
timestamp 1688980957
transform -1 0 421 0 1 0
box -260 1014 158 8958
use sky130_fd_io__tk_em1o_cdns_5595914180860  sky130_fd_io__tk_em1o_cdns_5595914180860_0
timestamp 1688980957
transform 0 -1 411 1 0 7019
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_0
timestamp 1688980957
transform 0 -1 409 1 0 9064
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_1
timestamp 1688980957
transform 0 -1 409 1 0 9624
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_2
timestamp 1688980957
transform 0 1 535 -1 0 10032
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_3
timestamp 1688980957
transform 0 1 535 -1 0 9451
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_4
timestamp 1688980957
transform 0 -1 411 1 0 8235
box 0 0 1 1
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_0
timestamp 1688980957
transform 0 -1 424 1 0 9101
box 15 13 285 14
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_1
timestamp 1688980957
transform 0 -1 424 1 0 9686
box 15 13 285 14
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_2
timestamp 1688980957
transform 0 1 520 -1 0 9966
box 15 13 285 14
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_3
timestamp 1688980957
transform 0 1 520 -1 0 9381
box 15 13 285 14
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1688980957
transform -1 0 397 0 1 9067
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1688980957
transform -1 0 397 0 -1 9665
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1688980957
transform 1 0 547 0 1 9632
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1688980957
transform 1 0 547 0 1 9047
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1688980957
transform 1 0 544 0 1 8772
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1688980957
transform 1 0 291 0 1 6332
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1688980957
transform 1 0 291 0 1 7674
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1688980957
transform -1 0 399 0 1 8908
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1688980957
transform 1 0 291 0 1 7566
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180857  sky130_fd_pr__via_l1m1__example_5595914180857_0
timestamp 1688980957
transform 1 0 468 0 1 5328
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_0
timestamp 1688980957
transform -1 0 397 0 1 9431
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_1
timestamp 1688980957
transform -1 0 397 0 -1 10099
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_2
timestamp 1688980957
transform 1 0 547 0 1 9994
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_3
timestamp 1688980957
transform 1 0 547 0 1 9442
box 0 0 1 1
<< labels >>
flabel metal1 s 479 5364 513 5398 0 FreeSans 200 0 0 0 RA
port 1 nsew
<< properties >>
string GDS_END 43499994
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43496546
<< end >>
