magic
tech sky130B
magscale 1 2
timestamp 1700463299
<< error_s >>
rect 4516 2259 4536 2460
rect 4544 2259 4564 2460
rect 4826 1748 4972 1760
rect 4872 1746 4972 1748
rect 4854 1718 5000 1732
rect 10014 738 10178 746
rect 10042 710 10206 718
rect 4796 -1122 4810 -790
rect 4792 -1172 4810 -1122
rect 4824 -1150 4838 -790
rect 4820 -1172 4838 -1150
rect 4792 -1428 4810 -1218
rect 4820 -1428 4838 -1218
rect 4792 -1678 4810 -1498
rect 4820 -1678 4838 -1498
rect 4792 -1766 4810 -1724
rect 4820 -1738 4838 -1724
rect 4798 -1938 4810 -1766
rect 4826 -1938 4838 -1738
<< metal1 >>
rect 8240 3576 8440 3584
rect 8240 3400 8252 3576
rect 8426 3400 8440 3576
rect 8240 3384 8440 3400
rect 4544 3254 4626 3264
rect 4542 3184 4552 3254
rect 4620 3184 4630 3254
rect 4544 3144 4626 3184
rect 4492 2944 4692 3144
rect 4544 1832 4626 2944
rect 4544 1830 4882 1832
rect 4534 1744 4544 1830
rect 4624 1748 4882 1830
rect 4624 1744 4634 1748
rect 4872 1746 4882 1748
rect 4962 1746 4972 1832
rect 13404 1746 13414 1922
rect 13588 1746 13598 1922
rect 4544 1736 4626 1744
rect 4600 600 5214 798
rect 4600 -2290 4810 600
rect 8474 300 8484 476
rect 8658 300 8668 476
rect 4600 -2322 5400 -2290
rect 4600 -2470 5568 -2322
rect 10296 -2470 10494 -958
rect 4600 -2488 10494 -2470
rect 5166 -2490 10494 -2488
rect 5366 -2676 10494 -2490
<< via1 >>
rect 8252 3400 8426 3576
rect 4552 3184 4620 3254
rect 4544 1744 4624 1830
rect 4882 1746 4962 1832
rect 13414 1746 13588 1922
rect 8484 300 8658 476
<< metal2 >>
rect 7984 3812 8090 3816
rect 7984 3746 10182 3812
rect 4490 3422 4690 3532
rect 7984 3422 8090 3746
rect 4490 3344 8090 3422
rect 8252 3576 8426 3586
rect 8252 3390 8426 3400
rect 4490 3332 4690 3344
rect 4552 3260 4620 3264
rect 4546 3254 5076 3260
rect 4546 3184 4552 3254
rect 4620 3184 5076 3254
rect 4546 3178 5076 3184
rect 4552 3174 4620 3178
rect 4888 2336 5088 2536
rect 4888 2002 5088 2202
rect 4544 1830 4624 1840
rect 4882 1836 4962 1842
rect 4544 1734 4624 1744
rect 4870 1832 4982 1836
rect 4870 1746 4882 1832
rect 4962 1746 4982 1832
rect 4870 168 4982 1746
rect 10100 1518 10182 3746
rect 13414 1922 13588 1932
rect 13414 1736 13588 1746
rect 9606 738 10178 828
rect 14730 512 14930 712
rect 8484 476 8658 486
rect 8484 290 8658 300
rect 9856 380 10172 478
rect 4870 70 5284 168
rect 5120 -752 5320 -552
rect 5118 -1084 5318 -884
rect 9856 -1100 9942 380
<< via2 >>
rect 8252 3400 8426 3576
rect 13414 1746 13588 1922
rect 8484 300 8658 476
<< metal3 >>
rect 8242 3576 8436 3581
rect 8242 3400 8252 3576
rect 8426 3574 8436 3576
rect 8426 3400 9842 3574
rect 8242 3395 8436 3400
rect 9668 1912 9840 3400
rect 13404 1922 13598 1927
rect 13404 1912 13414 1922
rect 9668 1746 13414 1912
rect 13588 1746 13598 1922
rect 9668 1741 13598 1746
rect 9668 1736 13584 1741
rect 8474 478 8668 481
rect 9668 478 9840 1736
rect 8474 476 9870 478
rect 8474 300 8484 476
rect 8658 302 9870 476
rect 8658 300 8668 302
rect 8474 295 8668 300
use 2-1MUX  x1
timestamp 1700463299
transform 1 0 5338 0 1 -3006
box -936 600 1824 2716
use 2-1MUX  x2
timestamp 1700463299
transform 1 0 5106 0 1 84
box -936 600 1824 2716
use 2-1MUX  x3
timestamp 1700463299
transform 1 0 10264 0 1 -1566
box -936 600 1824 2716
<< labels >>
flabel metal1 5166 -2490 5366 -2290 0 FreeSans 256 0 0 0 VSS
port 6 nsew
flabel metal1 4492 2944 4692 3144 0 FreeSans 256 0 0 0 S1
port 0 nsew
flabel metal1 8240 3384 8440 3584 0 FreeSans 256 0 0 0 VDD
port 5 nsew
flabel metal2 4490 3332 4690 3532 0 FreeSans 256 0 0 0 S2
port 8 nsew
flabel metal2 14730 512 14930 712 0 FreeSans 256 0 0 0 OUT
port 7 nsew
flabel metal2 5118 -1084 5318 -884 0 FreeSans 256 0 0 0 A
port 1 nsew
flabel metal2 4888 2002 5088 2202 0 FreeSans 256 0 0 0 C
port 3 nsew
flabel metal2 5120 -752 5320 -552 0 FreeSans 256 0 0 0 B
port 2 nsew
flabel metal2 4888 2336 5088 2536 0 FreeSans 256 0 0 0 D
port 4 nsew
<< end >>
