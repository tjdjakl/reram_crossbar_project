magic
tech sky130B
magscale 1 2
timestamp 1700625197
<< metal1 >>
rect 1462 2860 1662 2884
rect 1462 2700 1480 2860
rect 1640 2700 1662 2860
rect 1462 2684 1662 2700
rect 2508 2684 2708 2884
rect 4330 2720 4340 2880
rect 4500 2720 4510 2880
rect 4238 2382 4248 2492
rect 4384 2382 4394 2492
rect 1356 1794 1556 1846
rect 1356 1676 1384 1794
rect 1502 1676 1556 1794
rect 2066 1680 2076 1804
rect 2208 1680 2218 1804
rect 2408 1680 2418 1808
rect 2562 1680 2572 1808
rect 1356 1646 1556 1676
rect 4916 1642 5116 1842
rect 4242 1166 4252 1280
rect 4388 1166 4398 1280
rect 1460 850 1660 1050
rect 2148 828 2562 1116
rect 4147 1009 4437 1016
rect 4152 824 4346 1009
<< via1 >>
rect 1480 2700 1640 2860
rect 4340 2720 4500 2880
rect 4248 2382 4384 2492
rect 1384 1676 1502 1794
rect 2076 1680 2208 1804
rect 2418 1680 2562 1808
rect 4252 1166 4388 1280
<< metal2 >>
rect 4340 2880 4500 2890
rect 1480 2860 1640 2870
rect 4340 2710 4500 2720
rect 1480 2690 1640 2700
rect 4248 2492 4384 2502
rect 2076 2382 4248 2492
rect 4384 2382 4386 2492
rect 2076 1814 2206 2382
rect 4248 2372 4384 2382
rect 2076 1804 2208 1814
rect 1384 1794 1502 1804
rect 1384 1280 1502 1676
rect 2076 1670 2208 1680
rect 2418 1808 2562 1818
rect 2418 1670 2562 1680
rect 4252 1280 4388 1290
rect 1384 1166 4252 1280
rect 1384 1164 4388 1166
rect 4252 1156 4388 1164
<< via2 >>
rect 1480 2700 1640 2860
rect 4340 2720 4500 2880
rect 2418 1680 2562 1808
<< metal3 >>
rect 4330 2880 4510 2885
rect 1470 2860 1650 2865
rect 1470 2700 1480 2860
rect 1640 2700 1650 2860
rect 4330 2720 4340 2880
rect 4500 2720 4510 2880
rect 4330 2715 4510 2720
rect 1470 2695 1650 2700
rect 2408 1808 2572 1813
rect 2408 1680 2418 1808
rect 2562 1680 2572 1808
rect 2408 1675 2572 1680
rect 1180 1446 1380 1518
rect 2418 1446 2542 1675
rect 1180 1354 2542 1446
rect 1180 1318 1380 1354
<< via3 >>
rect 1480 2700 1640 2860
rect 4340 2720 4500 2880
<< metal4 >>
rect 4339 2880 4501 2881
rect 1520 2861 4340 2880
rect 1479 2860 4340 2861
rect 1479 2700 1480 2860
rect 1640 2720 4340 2860
rect 4500 2720 4501 2880
rect 1640 2719 4501 2720
rect 1640 2700 4460 2719
rect 1479 2699 1641 2700
use Buffer  x1
timestamp 1700618825
transform 1 0 544 0 1 -534
box 1858 1360 3698 3442
use TransmissionGate  x2
timestamp 1700624956
transform 1 0 4100 0 1 376
box 126 420 1016 2536
use Inverter  x3
timestamp 1700618825
transform 1 0 460 0 1 1270
box 896 -444 1780 1638
<< labels >>
flabel metal1 1356 1646 1556 1846 0 FreeSans 256 0 0 0 S
port 4 nsew
flabel metal3 1180 1318 1380 1518 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 1460 850 1660 1050 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 4916 1642 5116 1842 0 FreeSans 256 0 0 0 Vout
port 3 nsew
flabel metal1 2508 2684 2708 2884 0 FreeSans 256 0 0 0 VDD_25
port 5 nsew
flabel metal1 1462 2684 1662 2884 0 FreeSans 256 0 0 0 VDD_18
port 0 nsew
<< end >>
