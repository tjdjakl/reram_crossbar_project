magic
tech sky130B
magscale 1 2
timestamp 1700625197
<< metal1 >>
rect 27882 17688 28082 17888
rect 28928 17688 29128 17888
rect 29894 17700 29904 17856
rect 30046 17700 30056 17856
rect 27776 16650 27976 16850
rect 31336 16646 31536 16846
rect 27340 16510 27540 16522
rect 27340 16336 27476 16510
rect 27598 16336 27608 16510
rect 27340 16322 27540 16336
rect 27880 15854 28080 16054
rect 28930 15880 28940 16040
rect 29100 15880 29110 16040
rect 29904 15508 29914 15664
rect 30056 15508 30066 15664
rect 31336 14446 31536 14646
rect 27340 14310 27540 14322
rect 27340 14136 27472 14310
rect 27594 14136 27604 14310
rect 27340 14122 27540 14136
rect 28930 13680 28940 13840
rect 29100 13680 29110 13840
rect 29898 13304 29908 13460
rect 30050 13304 30060 13460
rect 31336 12246 31536 12446
rect 27340 12112 27540 12122
rect 27340 11938 27480 12112
rect 27602 11938 27612 12112
rect 27340 11922 27540 11938
rect 28930 11480 28940 11640
rect 29100 11480 29110 11640
rect 29896 11106 29906 11262
rect 30048 11106 30058 11262
rect 31336 10046 31536 10246
rect 27340 9910 27540 9922
rect 27340 9736 27476 9910
rect 27598 9736 27608 9910
rect 27340 9722 27540 9736
rect 28930 9280 28940 9440
rect 29100 9280 29110 9440
rect 29904 8898 29914 9054
rect 30056 8898 30066 9054
rect 31336 7846 31536 8046
rect 27340 7712 27540 7722
rect 27340 7538 27480 7712
rect 27602 7538 27612 7712
rect 27340 7522 27540 7538
rect 28930 7080 28940 7240
rect 29100 7080 29110 7240
rect 29906 6710 29916 6866
rect 30058 6710 30068 6866
rect 31336 5646 31536 5846
rect 27340 5508 27540 5522
rect 27340 5334 27480 5508
rect 27602 5334 27612 5508
rect 27340 5322 27540 5334
rect 28930 4880 28940 5040
rect 29100 4880 29110 5040
rect 29906 4504 29916 4660
rect 30058 4504 30068 4660
rect 31336 3446 31536 3646
rect 27360 3310 27560 3322
rect 27360 3136 27482 3310
rect 27604 3136 27614 3310
rect 27360 3122 27560 3136
rect 28930 2680 28940 2840
rect 29100 2680 29110 2840
rect 29910 2306 29920 2462
rect 30062 2306 30072 2462
rect 31336 1246 31536 1446
rect 27340 1110 27540 1122
rect 27340 936 27486 1110
rect 27608 936 27618 1110
rect 27340 922 27540 936
rect 28930 480 28940 640
rect 29100 480 29110 640
<< via1 >>
rect 29904 17700 30046 17856
rect 27476 16336 27598 16510
rect 28940 15880 29100 16040
rect 29914 15508 30056 15664
rect 27472 14136 27594 14310
rect 28940 13680 29100 13840
rect 29908 13304 30050 13460
rect 27480 11938 27602 12112
rect 28940 11480 29100 11640
rect 29906 11106 30048 11262
rect 27476 9736 27598 9910
rect 28940 9280 29100 9440
rect 29914 8898 30056 9054
rect 27480 7538 27602 7712
rect 28940 7080 29100 7240
rect 29916 6710 30058 6866
rect 27480 5334 27602 5508
rect 28940 4880 29100 5040
rect 29916 4504 30058 4660
rect 27482 3136 27604 3310
rect 28940 2680 29100 2840
rect 29920 2306 30062 2462
rect 27486 936 27608 1110
rect 28940 480 29100 640
<< metal2 >>
rect 29904 17856 30046 17866
rect 29904 17690 30046 17700
rect 27720 16726 27840 16800
rect 27476 16510 27598 16520
rect 27476 16326 27598 16336
rect 27472 14310 27594 14320
rect 27472 14126 27594 14136
rect 27480 12112 27602 12122
rect 27480 11928 27602 11938
rect 27476 9910 27598 9920
rect 27476 9726 27598 9736
rect 27480 7712 27602 7722
rect 27480 7528 27602 7538
rect 27480 5508 27602 5518
rect 27480 5324 27602 5334
rect 27482 3310 27604 3320
rect 27482 3126 27604 3136
rect 27720 1280 27842 16726
rect 28940 16040 29100 16050
rect 28940 15870 29100 15880
rect 29914 15664 30056 15674
rect 29914 15498 30056 15508
rect 28940 13840 29100 13850
rect 28940 13670 29100 13680
rect 29908 13460 30050 13470
rect 29908 13294 30050 13304
rect 28940 11640 29100 11650
rect 28940 11470 29100 11480
rect 29906 11262 30048 11272
rect 29906 11096 30048 11106
rect 28940 9440 29100 9450
rect 28940 9270 29100 9280
rect 29914 9054 30056 9064
rect 29914 8888 30056 8898
rect 28940 7240 29100 7250
rect 28940 7070 29100 7080
rect 29916 6866 30058 6876
rect 29916 6700 30058 6710
rect 28940 5040 29100 5050
rect 28940 4870 29100 4880
rect 29916 4660 30058 4670
rect 29916 4494 30058 4504
rect 28940 2840 29100 2850
rect 28940 2670 29100 2680
rect 29920 2462 30062 2472
rect 29920 2296 30062 2306
rect 27486 1110 27608 1120
rect 27486 926 27608 936
rect 28940 640 29100 650
rect 28940 470 29100 480
<< via2 >>
rect 29904 17700 30046 17856
rect 27476 16336 27598 16510
rect 27472 14136 27594 14310
rect 27480 11938 27602 12112
rect 27476 9736 27598 9910
rect 27480 7538 27602 7712
rect 27480 5334 27602 5508
rect 27482 3136 27604 3310
rect 28940 15880 29100 16040
rect 29914 15508 30056 15664
rect 28940 13680 29100 13840
rect 29908 13304 30050 13460
rect 28940 11480 29100 11640
rect 29906 11106 30048 11262
rect 28940 9280 29100 9440
rect 29914 8898 30056 9054
rect 28940 7080 29100 7240
rect 29916 6710 30058 6866
rect 28940 4880 29100 5040
rect 29916 4504 30058 4660
rect 28940 2680 29100 2840
rect 29920 2306 30062 2462
rect 27486 936 27608 1110
rect 28940 480 29100 640
<< metal3 >>
rect 29894 17856 30056 17861
rect 29894 17700 29904 17856
rect 30046 17764 30056 17856
rect 30046 17700 30062 17764
rect 29894 17695 30062 17700
rect 27466 16510 27608 16515
rect 27466 16336 27476 16510
rect 27598 16336 27608 16510
rect 27466 16331 27608 16336
rect 28930 16040 29110 16045
rect 28930 15880 28940 16040
rect 29100 15880 29720 16040
rect 28930 15875 29110 15880
rect 27462 14310 27604 14315
rect 27462 14136 27472 14310
rect 27594 14136 27604 14310
rect 27462 14131 27604 14136
rect 28930 13840 29110 13845
rect 29540 13840 29720 15880
rect 28930 13680 28940 13840
rect 29100 13680 29720 13840
rect 28930 13675 29110 13680
rect 27470 12112 27612 12117
rect 27470 11938 27480 12112
rect 27602 11938 27612 12112
rect 27470 11933 27612 11938
rect 28930 11640 29110 11645
rect 29540 11640 29720 13680
rect 29904 15669 30062 17695
rect 29904 15664 30066 15669
rect 29904 15508 29914 15664
rect 30056 15508 30066 15664
rect 29904 15503 30066 15508
rect 29904 13465 30062 15503
rect 29898 13460 30062 13465
rect 29898 13304 29908 13460
rect 30050 13304 30062 13460
rect 29898 13299 30062 13304
rect 28930 11480 28940 11640
rect 29100 11480 29720 11640
rect 28930 11475 29110 11480
rect 27466 9910 27608 9915
rect 27466 9736 27476 9910
rect 27598 9736 27608 9910
rect 27466 9731 27608 9736
rect 28930 9440 29110 9445
rect 29540 9440 29720 11480
rect 29904 11267 30062 13299
rect 29896 11262 30062 11267
rect 29896 11106 29906 11262
rect 30048 11106 30062 11262
rect 29896 11101 30062 11106
rect 28930 9280 28940 9440
rect 29100 9280 29720 9440
rect 28930 9275 29110 9280
rect 27470 7712 27612 7717
rect 27470 7538 27480 7712
rect 27602 7538 27612 7712
rect 27470 7533 27612 7538
rect 28930 7240 29110 7245
rect 29540 7240 29720 9280
rect 28930 7080 28940 7240
rect 29100 7080 29720 7240
rect 28930 7075 29110 7080
rect 27470 5508 27612 5513
rect 27470 5334 27480 5508
rect 27602 5334 27612 5508
rect 27470 5329 27612 5334
rect 28930 5040 29110 5045
rect 29540 5040 29720 7080
rect 28930 4880 28940 5040
rect 29100 4880 29720 5040
rect 28930 4875 29110 4880
rect 27472 3310 27614 3315
rect 27472 3136 27482 3310
rect 27604 3136 27614 3310
rect 27472 3131 27614 3136
rect 28930 2840 29110 2845
rect 29540 2840 29720 4880
rect 28930 2680 28940 2840
rect 29100 2680 29720 2840
rect 28930 2675 29110 2680
rect 27476 1110 27618 1115
rect 27476 936 27486 1110
rect 27608 936 27618 1110
rect 27476 931 27618 936
rect 28930 640 29110 645
rect 29540 640 29720 2680
rect 29904 9059 30062 11101
rect 29904 9054 30066 9059
rect 29904 8898 29914 9054
rect 30056 8898 30066 9054
rect 29904 8893 30066 8898
rect 29904 6871 30062 8893
rect 29904 6866 30068 6871
rect 29904 6710 29916 6866
rect 30058 6710 30068 6866
rect 29904 6705 30068 6710
rect 29904 4665 30062 6705
rect 29904 4660 30068 4665
rect 29904 4504 29916 4660
rect 30058 4504 30068 4660
rect 29904 4499 30068 4504
rect 29904 2467 30062 4499
rect 29904 2462 30072 2467
rect 29904 2386 29920 2462
rect 29910 2306 29920 2386
rect 30062 2306 30072 2462
rect 29910 2301 30072 2306
rect 28930 480 28940 640
rect 29100 480 29720 640
rect 28930 475 29110 480
<< metal4 >>
rect 30760 2380 30920 17820
use 1LineSelectInput  x1
timestamp 1700625197
transform 1 0 26420 0 1 15004
box 1180 796 5116 2912
use 1LineSelectInput  x2
timestamp 1700625197
transform 1 0 26420 0 1 12804
box 1180 796 5116 2912
use 1LineSelectInput  x3
timestamp 1700625197
transform 1 0 26420 0 1 10604
box 1180 796 5116 2912
use 1LineSelectInput  x4
timestamp 1700625197
transform 1 0 26420 0 1 8404
box 1180 796 5116 2912
use 1LineSelectInput  x5
timestamp 1700625197
transform 1 0 26420 0 1 6204
box 1180 796 5116 2912
use 1LineSelectInput  x6
timestamp 1700625197
transform 1 0 26420 0 1 4004
box 1180 796 5116 2912
use 1LineSelectInput  x7
timestamp 1700625197
transform 1 0 26420 0 1 1804
box 1180 796 5116 2912
use 1LineSelectInput  x8
timestamp 1700625197
transform 1 0 26420 0 1 -396
box 1180 796 5116 2912
<< labels >>
flabel metal1 27776 16650 27976 16850 0 FreeSans 256 0 0 0 S
port 11 nsew
flabel metal1 31336 16646 31536 16846 0 FreeSans 256 0 0 0 SL_IN1
port 19 nsew
flabel metal1 31336 14446 31536 14646 0 FreeSans 256 0 0 0 SL_IN2
port 18 nsew
flabel metal1 31336 12246 31536 12446 0 FreeSans 256 0 0 0 SL_IN3
port 17 nsew
flabel metal1 31336 10046 31536 10246 0 FreeSans 256 0 0 0 SL_IN4
port 16 nsew
flabel metal1 31336 7846 31536 8046 0 FreeSans 256 0 0 0 SL_IN5
port 15 nsew
flabel metal1 31336 5646 31536 5846 0 FreeSans 256 0 0 0 SL_IN6
port 14 nsew
flabel metal1 31336 3446 31536 3646 0 FreeSans 256 0 0 0 SL_IN7
port 13 nsew
flabel metal1 31336 1246 31536 1446 0 FreeSans 256 0 0 0 SL_IN8
port 12 nsew
flabel metal1 27880 15854 28080 16054 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 27340 922 27540 1122 0 FreeSans 256 0 0 0 SL_LA_IN8
port 2 nsew
flabel metal1 27360 3122 27560 3322 0 FreeSans 256 0 0 0 SL_LA_IN7
port 3 nsew
flabel metal1 27340 5322 27540 5522 0 FreeSans 256 0 0 0 SL_LA_IN6
port 4 nsew
flabel metal1 27340 7522 27540 7722 0 FreeSans 256 0 0 0 SL_LA_IN5
port 5 nsew
flabel metal1 27340 9722 27540 9922 0 FreeSans 256 0 0 0 SL_LA_IN4
port 6 nsew
flabel metal1 27340 11922 27540 12122 0 FreeSans 256 0 0 0 SL_LA_IN3
port 7 nsew
flabel metal1 27340 14122 27540 14322 0 FreeSans 256 0 0 0 SL_LA_IN2
port 9 nsew
flabel metal1 27340 16322 27540 16522 0 FreeSans 256 0 0 0 SL_LA_IN1
port 10 nsew
flabel metal1 28928 17688 29128 17888 0 FreeSans 256 0 0 0 VDD25
port 0 nsew
flabel metal1 27882 17688 28082 17888 0 FreeSans 256 0 0 0 VDD18
port 20 nsew
<< end >>
