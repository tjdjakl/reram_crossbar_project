magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< obsli1 >>
rect 48 204 14951 39556
<< metal1 >>
rect 5242 0 5540 34
<< obsm1 >>
rect 24 90 14957 39568
rect 24 0 5186 90
rect 5596 0 14957 90
<< metal2 >>
rect 100 0 4099 297
rect 6888 0 8888 65
rect 10943 0 14940 732
<< obsm2 >>
rect 100 788 14940 38886
rect 100 353 10887 788
rect 4155 121 10887 353
rect 4155 0 6832 121
rect 8944 0 10887 121
<< metal3 >>
rect 1009 11667 1011 11669
rect 13489 11667 13491 11669
rect 100 0 4900 11064
rect 5200 0 7376 4044
rect 7676 0 9851 4580
rect 10151 0 14940 11064
<< obsm3 >>
rect 100 11749 14940 37903
rect 100 11587 929 11749
rect 1091 11587 13409 11749
rect 13571 11587 14940 11749
rect 100 11144 14940 11587
rect 4980 4660 10071 11144
rect 4980 4124 7596 4660
rect 4980 3558 5120 4124
rect 7456 3558 7596 4124
rect 9931 3558 10071 4660
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 15000 10947
rect 0 10225 254 10821
rect 0 9929 254 10165
rect 0 9273 254 9869
rect 14746 10225 15000 10821
rect 14746 9929 15000 10165
rect 14746 9273 15000 9869
rect 0 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< obsm4 >>
rect 334 34677 14666 39600
rect 193 18680 14807 34677
rect 334 13527 14666 18680
rect 193 13387 14807 13527
rect 334 12337 14666 13387
rect 193 12217 14807 12337
rect 334 11167 14666 12217
rect 193 11027 14807 11167
rect 334 9293 14666 10801
rect 193 8927 14807 9067
rect 334 7837 14666 8927
rect 193 7717 14807 7837
rect 334 6867 14666 7717
rect 193 6747 14807 6867
rect 334 5897 14666 6747
rect 193 5777 14807 5897
rect 334 4687 14666 5777
rect 193 4567 14807 4687
rect 334 3477 14666 4567
rect 193 3357 14807 3477
rect 273 2507 14727 3357
rect 193 2387 14807 2507
rect 334 1297 14666 2387
rect 193 1177 14807 1297
rect 334 7 14666 1177
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 2054 33433 2082 33461
rect 0 13607 254 18597
rect 0 12437 254 13287
rect 0 11267 254 12117
rect 0 9147 254 10947
rect 0 7937 254 8827
rect 0 6968 254 7617
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 11267 15000 12117
rect 14746 9147 15000 10947
rect 14746 7937 15000 8827
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 0 4787 254 5677
rect 0 3577 254 4467
rect 14746 5997 15000 6647
rect 14746 4787 15000 5677
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 0 27 254 1077
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 574 34437 14426 39600
rect 0 33781 15000 34437
rect 0 33113 1734 33781
rect 2402 33113 15000 33781
rect 0 18917 15000 33113
rect 574 6968 14426 18917
rect 0 6967 15000 6968
rect 574 3257 14426 6967
rect 513 2607 14487 3257
rect 574 27 14426 2607
<< labels >>
rlabel metal3 s 13489 11667 13491 11669 6 PADISOR
port 1 nsew
rlabel metal3 s 1009 11667 1011 11669 6 PADISOL
port 2 nsew
rlabel metal4 s 0 4767 254 5697 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal4 s 0 34757 254 39600 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 9147 15000 9213 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 10881 15000 10947 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 6947 254 7637 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 11247 254 12137 6 VSSIO_Q
port 5 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 VSSIO_Q
port 5 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 5 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 5 nsew ground bidirectional
rlabel metal4 s 0 7 254 1097 6 VCCHIB
port 6 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 VCCHIB
port 6 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 6 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 6 nsew power bidirectional
rlabel metal4 s 0 1377 254 2307 6 VCCD
port 7 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 7 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 7 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 7 nsew power bidirectional
rlabel metal4 s 0 2587 193 3277 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 0 3557 254 4487 6 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 6 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 6 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 6 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 0 5977 254 6667 6 VSWITCH
port 10 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 10 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 10 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 10 nsew power bidirectional
rlabel metal4 s 0 12417 254 13307 6 VDDIO_Q
port 11 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 6 VDDIO_Q
port 11 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 11 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 11 nsew power bidirectional
rlabel metal4 s 0 10225 254 10821 6 AMUXBUS_A
port 12 nsew signal bidirectional
rlabel metal4 s 14746 10225 15000 10821 6 AMUXBUS_A
port 12 nsew signal bidirectional
rlabel metal4 s 0 9273 254 9869 6 AMUXBUS_B
port 13 nsew signal bidirectional
rlabel metal4 s 14746 9273 15000 9869 6 AMUXBUS_B
port 13 nsew signal bidirectional
rlabel metal4 s 0 7917 254 8847 6 VSSD
port 14 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 14 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 14 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 14 nsew ground bidirectional
rlabel metal5 s 2054 33433 2082 33461 6 G_PAD
port 15 nsew signal bidirectional
rlabel metal2 s 100 0 4099 297 6 SRC_BDY_LVC1
port 16 nsew ground bidirectional
rlabel metal2 s 10943 0 14940 732 6 SRC_BDY_LVC2
port 17 nsew ground bidirectional
rlabel metal2 s 6888 0 8888 65 6 BDY2_B2B
port 18 nsew ground bidirectional
rlabel metal3 s 7676 0 9851 4580 6 DRN_LVC2
port 19 nsew power bidirectional
rlabel metal3 s 5200 0 7376 4044 6 DRN_LVC1
port 20 nsew power bidirectional
rlabel metal3 s 10151 0 14940 11064 6 G_CORE
port 21 nsew ground bidirectional
rlabel metal3 s 100 0 4900 11064 6 G_CORE
port 21 nsew ground bidirectional
rlabel metal1 s 5242 0 5540 34 6 OGC_LVC
port 22 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 19149052
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 15530004
<< end >>
