magic
tech sky130B
timestamp 1688980957
<< properties >>
string GDS_END 3163080
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3162756
<< end >>
