magic
tech sky130B
magscale 1 2
timestamp 1700640585
<< metal1 >>
rect 58616 62742 58816 62942
rect 69890 60551 70090 60751
rect 57552 59058 57752 59258
rect 66980 59150 67180 59350
rect 57310 58620 57320 58780
rect 57480 58620 57490 58780
rect 58950 58735 59150 58935
rect 69889 48552 70089 48752
rect 57310 46620 57320 46780
rect 57480 46620 57490 46780
rect 69890 36552 70090 36752
rect 57310 34620 57320 34780
rect 57480 34620 57490 34780
rect 69890 24552 70090 24752
rect 57310 22620 57320 22780
rect 57480 22620 57490 22780
rect 32179 14776 32379 14976
rect 46052 14708 46252 14908
rect 44610 13680 44620 13840
rect 44780 13680 44790 13840
rect 48596 13343 48796 13543
rect 32180 12576 32380 12776
rect 69890 12551 70090 12751
rect 44610 11480 44620 11640
rect 44780 11480 44790 11640
rect 48596 11142 48796 11342
rect 57310 10620 57320 10780
rect 57480 10620 57490 10780
rect 32180 10376 32380 10576
rect 44610 9280 44620 9440
rect 44780 9280 44790 9440
rect 48596 8942 48796 9142
rect 32181 8176 32381 8376
rect 44610 7080 44620 7240
rect 44780 7080 44790 7240
rect 48596 6742 48796 6942
rect 32180 5976 32380 6176
rect 44610 4880 44620 5040
rect 44780 4880 44790 5040
rect 48596 4542 48796 4742
rect 32180 3776 32380 3976
rect 44610 2680 44620 2840
rect 44780 2680 44790 2840
rect 48596 2342 48796 2542
rect 32180 1576 32380 1776
rect 44610 480 44620 640
rect 44780 480 44790 640
rect 69890 552 70090 752
rect 48575 142 48775 342
rect 32181 -624 32381 -424
rect 45188 -672 45388 -472
rect 57310 -1380 57320 -1220
rect 57480 -1380 57490 -1220
rect 44610 -1720 44620 -1560
rect 44780 -1720 44790 -1560
rect 48160 -1730 48360 -1530
rect 32393 -2016 32593 -1816
rect 48596 -2058 48796 -1858
rect 30432 -2389 30632 -2189
rect 47012 -2526 47212 -2326
rect 30420 -2855 30620 -2655
rect 30431 -3502 30631 -3302
rect 32392 -3912 32592 -3712
rect 30486 -4531 30686 -4331
rect 30392 -4922 30592 -4722
rect 30380 -5568 30580 -5368
rect 30392 -6034 30592 -5834
rect 30484 -6364 30684 -6164
rect 32835 -7780 33035 -7580
rect 34484 -7759 34494 -7619
rect 34654 -7759 34664 -7619
rect 32836 -10180 33036 -9980
rect 34483 -10160 34493 -10020
rect 34653 -10160 34663 -10020
rect 69890 -11448 70090 -11248
rect 32836 -12580 33036 -12380
rect 34479 -12557 34489 -12417
rect 34649 -12557 34659 -12417
rect 57310 -13380 57320 -13220
rect 57480 -13380 57490 -13220
rect 32836 -14980 33036 -14780
rect 34483 -14954 34493 -14814
rect 34653 -14954 34663 -14814
rect 32836 -17380 33036 -17180
rect 34488 -17347 34498 -17207
rect 34658 -17347 34668 -17207
rect 32836 -19780 33036 -19580
rect 34486 -19749 34496 -19609
rect 34656 -19749 34666 -19609
rect 32836 -22180 33036 -21980
rect 34488 -22151 34498 -22011
rect 34658 -22151 34668 -22011
rect 69890 -23448 70090 -23248
rect 32836 -24580 33036 -24380
rect 34490 -24560 34500 -24420
rect 34660 -24560 34670 -24420
rect 38140 -24980 38340 -24780
rect 57310 -25380 57320 -25220
rect 57480 -25380 57490 -25220
<< via1 >>
rect 57320 58620 57480 58780
rect 57320 46620 57480 46780
rect 57320 34620 57480 34780
rect 57320 22620 57480 22780
rect 44620 13680 44780 13840
rect 44620 11480 44780 11640
rect 57320 10620 57480 10780
rect 44620 9280 44780 9440
rect 44620 7080 44780 7240
rect 44620 4880 44780 5040
rect 44620 2680 44780 2840
rect 44620 480 44780 640
rect 57320 -1380 57480 -1220
rect 44620 -1720 44780 -1560
rect 34494 -7759 34654 -7619
rect 34493 -10160 34653 -10020
rect 34489 -12557 34649 -12417
rect 57320 -13380 57480 -13220
rect 34493 -14954 34653 -14814
rect 34498 -17347 34658 -17207
rect 34496 -19749 34656 -19609
rect 34498 -22151 34658 -22011
rect 34500 -24560 34660 -24420
rect 57320 -25380 57480 -25220
<< metal2 >>
rect 57320 58780 57480 58790
rect 38200 58620 57320 58780
rect 37714 14908 37854 14918
rect 37714 14796 37854 14806
rect 38200 13520 38360 58620
rect 57320 58610 57480 58620
rect 57320 46780 57480 46790
rect 38200 13350 38360 13360
rect 38880 46620 57320 46780
rect 37714 12708 37854 12718
rect 37714 12596 37854 12606
rect 38880 11320 39040 46620
rect 57320 46610 57480 46620
rect 57320 34780 57480 34790
rect 38880 11170 39040 11180
rect 39580 34620 57320 34780
rect 37714 10508 37854 10518
rect 37714 10396 37854 10406
rect 39580 9180 39740 34620
rect 57320 34610 57480 34620
rect 57320 22780 57480 22790
rect 39580 9010 39740 9020
rect 40280 22620 57320 22780
rect 37714 8308 37854 8318
rect 37714 8196 37854 8206
rect 40280 7080 40440 22620
rect 57320 22610 57480 22620
rect 44620 13840 44780 13850
rect 44620 13670 44780 13680
rect 44620 11640 44780 11650
rect 44620 11470 44780 11480
rect 57320 10780 57480 10790
rect 54760 10620 57320 10780
rect 54760 10610 57480 10620
rect 54760 10600 57400 10610
rect 44620 9440 44780 9450
rect 44620 9270 44780 9280
rect 44620 7240 44780 7250
rect 44620 7070 44780 7080
rect 40280 6910 40440 6920
rect 37714 6108 37854 6118
rect 37714 5996 37854 6006
rect 44620 5040 44780 5050
rect 44620 4870 44780 4880
rect 37714 3908 37854 3918
rect 37714 3796 37854 3806
rect 44620 2840 44780 2850
rect 44620 2670 44780 2680
rect 37714 1708 37854 1718
rect 37714 1596 37854 1606
rect 44620 640 44780 650
rect 44620 470 44780 480
rect 32180 -203 32380 -3
rect 37714 -492 37854 -482
rect 37714 -604 37854 -594
rect 32180 -1044 32380 -844
rect 44620 -1560 44780 -1550
rect 44620 -1730 44780 -1720
rect 40960 -4960 41120 -4950
rect 54760 -4960 55040 10600
rect 57320 -1220 57480 -1210
rect 41120 -5120 55040 -4960
rect 55500 -1380 57320 -1220
rect 40960 -5130 41120 -5120
rect 41660 -5380 41820 -5370
rect 55500 -5380 55740 -1380
rect 57320 -1390 57480 -1380
rect 41820 -5540 55740 -5380
rect 41660 -5550 41820 -5540
rect 42360 -5720 42520 -5710
rect 42520 -5880 44560 -5720
rect 42360 -5890 42520 -5880
rect 43060 -6140 43220 -6130
rect 43220 -6300 44000 -6140
rect 43060 -6310 43220 -6300
rect 34494 -7619 34654 -7609
rect 34654 -7627 36425 -7626
rect 34654 -7629 37771 -7627
rect 34654 -7759 37772 -7629
rect 34494 -7761 37772 -7759
rect 34494 -7763 36425 -7761
rect 34494 -7769 34654 -7763
rect 37602 -8413 37772 -7761
rect 37602 -8529 38085 -8413
rect 34493 -10014 34653 -10010
rect 36514 -10013 37798 -10011
rect 36514 -10014 37845 -10013
rect 34493 -10020 37845 -10014
rect 34653 -10148 37845 -10020
rect 34493 -10170 34653 -10160
rect 37678 -10716 37845 -10148
rect 37676 -10830 38131 -10716
rect 34489 -12417 34649 -12407
rect 36334 -12413 37652 -12412
rect 36334 -12421 37812 -12413
rect 34649 -12555 37812 -12421
rect 34489 -12567 34649 -12557
rect 37616 -12997 37812 -12555
rect 37616 -13118 38090 -12997
rect 34493 -14814 34653 -14804
rect 36314 -14814 37782 -14812
rect 36314 -14824 37784 -14814
rect 34653 -14954 37784 -14824
rect 34493 -14958 37784 -14954
rect 34493 -14964 34653 -14958
rect 37642 -15311 37784 -14958
rect 37642 -15428 38120 -15311
rect 37644 -15436 38120 -15428
rect 34498 -17207 34658 -17197
rect 36414 -17214 37733 -17212
rect 36414 -17220 37734 -17214
rect 34658 -17347 37734 -17220
rect 34498 -17354 37734 -17347
rect 34498 -17357 34658 -17354
rect 36414 -17355 37734 -17354
rect 37518 -17597 37734 -17355
rect 37518 -17720 38100 -17597
rect 34496 -19609 34656 -19599
rect 36334 -19620 37847 -19604
rect 34656 -19749 37847 -19620
rect 34496 -19753 37847 -19749
rect 34496 -19754 37664 -19753
rect 34496 -19759 34656 -19754
rect 37697 -19919 37847 -19753
rect 37697 -20031 38131 -19919
rect 34498 -22011 34658 -22001
rect 36394 -22024 37728 -22018
rect 34658 -22151 37728 -22024
rect 34498 -22158 37728 -22151
rect 34498 -22161 34658 -22158
rect 37554 -22193 37728 -22158
rect 37554 -22317 38113 -22193
rect 34500 -24420 34660 -24410
rect 36354 -24450 38088 -24433
rect 34660 -24560 38088 -24450
rect 34500 -24570 38141 -24560
rect 34572 -24584 38141 -24570
rect 36354 -24590 38141 -24584
rect 43840 -25220 44000 -6300
rect 44360 -13220 44560 -5880
rect 57320 -13220 57480 -13210
rect 44360 -13380 57320 -13220
rect 57320 -13390 57480 -13380
rect 57320 -25220 57480 -25210
rect 43840 -25380 57320 -25220
rect 57320 -25390 57480 -25380
<< via2 >>
rect 37714 14806 37854 14908
rect 38200 13360 38360 13520
rect 37714 12606 37854 12708
rect 38880 11180 39040 11320
rect 37714 10406 37854 10508
rect 39580 9020 39740 9180
rect 37714 8206 37854 8308
rect 44620 13680 44780 13840
rect 44620 11480 44780 11640
rect 44620 9280 44780 9440
rect 40280 6920 40440 7080
rect 44620 7080 44780 7240
rect 37714 6006 37854 6108
rect 44620 4880 44780 5040
rect 37714 3806 37854 3908
rect 44620 2680 44780 2840
rect 37714 1606 37854 1708
rect 44620 480 44780 640
rect 37714 -594 37854 -492
rect 44620 -1720 44780 -1560
rect 40960 -5120 41120 -4960
rect 41660 -5540 41820 -5380
rect 42360 -5880 42520 -5720
rect 43060 -6300 43220 -6140
<< metal3 >>
rect 37704 14908 37864 14913
rect 37704 14806 37714 14908
rect 37854 14806 37864 14908
rect 37704 14801 37864 14806
rect 44610 13840 44790 13845
rect 38200 13680 44620 13840
rect 44780 13680 44790 13840
rect 38200 13525 38360 13680
rect 44610 13675 44790 13680
rect 38190 13520 38370 13525
rect 38190 13360 38200 13520
rect 38360 13360 38370 13520
rect 38190 13355 38370 13360
rect 37704 12708 37864 12713
rect 37704 12606 37714 12708
rect 37854 12606 37864 12708
rect 37704 12601 37864 12606
rect 37704 10508 37864 10513
rect 37704 10406 37714 10508
rect 37854 10406 37864 10508
rect 37704 10401 37864 10406
rect 37704 8308 37864 8313
rect 37704 8206 37714 8308
rect 37854 8206 37864 8308
rect 37704 8201 37864 8206
rect 37704 6108 37864 6113
rect 37704 6006 37714 6108
rect 37854 6006 37864 6108
rect 37704 6001 37864 6006
rect 37704 3908 37864 3913
rect 37704 3806 37714 3908
rect 37854 3806 37864 3908
rect 37704 3801 37864 3806
rect 37704 1708 37864 1713
rect 37704 1606 37714 1708
rect 37854 1606 37864 1708
rect 37704 1601 37864 1606
rect 37704 -492 37864 -487
rect 37704 -594 37714 -492
rect 37854 -594 37864 -492
rect 37704 -599 37864 -594
rect 38200 -6740 38360 13355
rect 44610 11640 44790 11645
rect 38880 11480 44620 11640
rect 44780 11480 44790 11640
rect 38880 11475 44790 11480
rect 38880 11460 44700 11475
rect 38880 11345 39040 11460
rect 38870 11320 39050 11345
rect 38870 11180 38880 11320
rect 39040 11180 39050 11320
rect 38870 11175 39050 11180
rect 38450 -6820 38460 -6708
rect 38618 -6820 38628 -6708
rect 38880 -6720 39040 11175
rect 44610 9440 44790 9445
rect 39580 9280 44620 9440
rect 44780 9280 44790 9440
rect 39580 9185 39740 9280
rect 44610 9275 44790 9280
rect 39570 9180 39750 9185
rect 39570 9020 39580 9180
rect 39740 9020 39750 9180
rect 39570 9015 39750 9020
rect 39144 -6820 39154 -6708
rect 39312 -6820 39322 -6708
rect 39580 -6800 39740 9015
rect 44610 7240 44790 7245
rect 40280 7085 44620 7240
rect 40270 7080 44620 7085
rect 44780 7080 44790 7240
rect 40270 6920 40280 7080
rect 40440 6920 40450 7080
rect 44610 7075 44790 7080
rect 40270 6915 40450 6920
rect 39842 -6820 39852 -6708
rect 40010 -6820 40020 -6708
rect 40280 -6800 40440 6915
rect 44610 5040 44790 5045
rect 40960 4880 44620 5040
rect 44780 4880 44790 5040
rect 40960 -4955 41120 4880
rect 44610 4875 44790 4880
rect 44610 2840 44790 2845
rect 41660 2680 44620 2840
rect 44780 2680 44790 2840
rect 40950 -4960 41130 -4955
rect 40950 -5120 40960 -4960
rect 41120 -5120 41130 -4960
rect 40950 -5125 41130 -5120
rect 40536 -6820 40546 -6708
rect 40704 -6820 40714 -6708
rect 40960 -6760 41120 -5125
rect 41660 -5375 41820 2680
rect 44610 2675 44790 2680
rect 44610 640 44790 645
rect 42360 480 44620 640
rect 44780 480 44790 640
rect 41650 -5380 41830 -5375
rect 41650 -5540 41660 -5380
rect 41820 -5540 41830 -5380
rect 41650 -5545 41830 -5540
rect 41226 -6820 41236 -6708
rect 41394 -6820 41404 -6708
rect 41660 -6740 41820 -5545
rect 42360 -5715 42520 480
rect 44610 475 44790 480
rect 44610 -1560 44790 -1555
rect 43060 -1720 44620 -1560
rect 44780 -1720 44790 -1560
rect 42350 -5720 42530 -5715
rect 42350 -5880 42360 -5720
rect 42520 -5880 42530 -5720
rect 42350 -5885 42530 -5880
rect 41920 -6820 41930 -6708
rect 42088 -6820 42098 -6708
rect 42360 -6820 42520 -5885
rect 43060 -6135 43220 -1720
rect 44610 -1725 44790 -1720
rect 43050 -6140 43230 -6135
rect 43050 -6300 43060 -6140
rect 43220 -6300 43230 -6140
rect 43050 -6305 43230 -6300
rect 42618 -6820 42628 -6708
rect 42786 -6820 42796 -6708
rect 43060 -6780 43220 -6305
rect 43312 -6820 43322 -6708
rect 43480 -6820 43490 -6708
<< via3 >>
rect 37714 14806 37854 14908
rect 37714 12606 37854 12708
rect 37714 10406 37854 10508
rect 37714 8206 37854 8308
rect 37714 6006 37854 6108
rect 37714 3806 37854 3908
rect 37714 1606 37854 1708
rect 37714 -594 37854 -492
rect 38460 -6820 38618 -6708
rect 39154 -6820 39312 -6708
rect 39852 -6820 40010 -6708
rect 40546 -6820 40704 -6708
rect 41236 -6820 41394 -6708
rect 41930 -6820 42088 -6708
rect 42628 -6820 42786 -6708
rect 43322 -6820 43480 -6708
<< metal4 >>
rect 37700 14908 43520 14920
rect 37700 14806 37714 14908
rect 37854 14806 43520 14908
rect 37700 14800 43520 14806
rect 37720 12709 42800 12720
rect 37713 12708 42800 12709
rect 37713 12606 37714 12708
rect 37854 12606 42800 12708
rect 37713 12605 42800 12606
rect 37720 12600 42800 12605
rect 37720 10509 42080 10520
rect 37713 10508 42080 10509
rect 37713 10406 37714 10508
rect 37854 10406 42080 10508
rect 37713 10405 42080 10406
rect 37720 10400 42080 10405
rect 37720 8309 41400 8320
rect 37713 8308 41400 8309
rect 37713 8206 37714 8308
rect 37854 8206 41400 8308
rect 37713 8205 41400 8206
rect 37720 8200 41400 8205
rect 37740 6109 40700 6120
rect 37713 6108 40700 6109
rect 37713 6006 37714 6108
rect 37854 6006 40700 6108
rect 37713 6005 40700 6006
rect 37740 6000 40700 6005
rect 37760 3909 40020 3920
rect 37713 3908 40020 3909
rect 37713 3806 37714 3908
rect 37854 3806 40020 3908
rect 37713 3805 40020 3806
rect 37760 3800 40020 3805
rect 37740 1709 39320 1720
rect 37713 1708 39320 1709
rect 37713 1606 37714 1708
rect 37854 1606 39320 1708
rect 37713 1605 39320 1606
rect 37740 1600 39320 1605
rect 37700 -492 38620 -480
rect 37700 -594 37714 -492
rect 37854 -594 38620 -492
rect 37700 -600 38620 -594
rect 38460 -6707 38620 -600
rect 39160 -6707 39320 1600
rect 39860 -6707 40020 3800
rect 38459 -6708 38620 -6707
rect 38459 -6820 38460 -6708
rect 38618 -6780 38620 -6708
rect 39153 -6708 39320 -6707
rect 38618 -6820 38619 -6780
rect 38459 -6821 38619 -6820
rect 39153 -6820 39154 -6708
rect 39312 -6800 39320 -6708
rect 39851 -6708 40020 -6707
rect 39312 -6820 39313 -6800
rect 39153 -6821 39313 -6820
rect 39851 -6820 39852 -6708
rect 40010 -6740 40020 -6708
rect 40540 -6707 40700 6000
rect 41240 -6707 41400 8200
rect 40540 -6708 40705 -6707
rect 40540 -6720 40546 -6708
rect 40010 -6820 40011 -6740
rect 39851 -6821 40011 -6820
rect 40545 -6820 40546 -6720
rect 40704 -6820 40705 -6708
rect 40545 -6821 40705 -6820
rect 41235 -6708 41400 -6707
rect 41235 -6820 41236 -6708
rect 41394 -6720 41400 -6708
rect 41920 -6707 42080 10400
rect 42640 -6707 42800 12600
rect 43340 12540 43520 14800
rect 43340 -6707 43500 12540
rect 41920 -6708 42089 -6707
rect 41920 -6720 41930 -6708
rect 41394 -6820 41395 -6720
rect 41235 -6821 41395 -6820
rect 41929 -6820 41930 -6720
rect 42088 -6820 42089 -6708
rect 41929 -6821 42089 -6820
rect 42627 -6708 42800 -6707
rect 42627 -6820 42628 -6708
rect 42786 -6740 42800 -6708
rect 43321 -6708 43500 -6707
rect 42786 -6820 42787 -6740
rect 42627 -6821 42787 -6820
rect 43321 -6820 43322 -6708
rect 43480 -6740 43500 -6708
rect 43480 -6820 43481 -6740
rect 43321 -6821 43481 -6820
use 64T64R  x1
timestamp 1700618825
transform 1 0 24980 0 1 -23036
box 13020 -1964 18566 16364
use 8LineSelectInput  x2
timestamp 1700625197
transform -1 0 76136 0 1 -2980
box 27340 400 31536 17916
use 8LineWordInput  x3
timestamp 1700640585
transform 1 0 33036 0 1 -27200
box -2656 1800 1640 22896
use 8LineBitInput  x4
timestamp 1700640585
transform 1 0 -980 0 -1 19196
box 31400 3400 38864 23116
use 8LineSelectOutput02  x5
timestamp 1700618825
transform 1 0 -33000 0 1 -25800
box 90200 400 103090 96282
<< labels >>
flabel metal1 32181 -624 32381 -424 0 FreeSans 256 0 0 0 {la_data_in\[0\]}
port 9 nsew
flabel metal1 32180 1576 32380 1776 0 FreeSans 256 0 0 0 {la_data_in\[1\]}
port 10 nsew
flabel metal1 32180 3776 32380 3976 0 FreeSans 256 0 0 0 {la_data_in\[2\]}
port 11 nsew
flabel metal1 32180 5976 32380 6176 0 FreeSans 256 0 0 0 {la_data_in\[3\]}
port 12 nsew
flabel metal1 32181 8176 32381 8376 0 FreeSans 256 0 0 0 {la_data_in\[4\]}
port 13 nsew
flabel metal1 32180 10376 32380 10576 0 FreeSans 256 0 0 0 {la_data_in\[5\]}
port 15 nsew
flabel metal1 32180 12576 32380 12776 0 FreeSans 256 0 0 0 {la_data_in\[6\]}
port 16 nsew
flabel metal1 32179 14776 32379 14976 0 FreeSans 256 0 0 0 {la_data_in\[7\]}
port 17 nsew
flabel metal2 32180 -203 32380 -3 0 FreeSans 256 0 0 0 v02B
port 34 nsew
flabel metal1 30420 -2855 30620 -2655 0 FreeSans 256 0 0 0 {la_data_in\[24\]B}
port 27 nsew
flabel metal1 30431 -3502 30631 -3302 0 FreeSans 256 0 0 0 v25B
port 32 nsew
flabel metal1 30432 -2389 30632 -2189 0 FreeSans 256 0 0 0 v3B
port 33 nsew
flabel metal1 32392 -3912 32592 -3712 0 FreeSans 256 0 0 0 vddB
port 37 nsew
flabel metal1 32393 -2016 32593 -1816 0 FreeSans 256 0 0 0 vssB
port 38 nsew
flabel metal1 30484 -6364 30684 -6164 0 FreeSans 256 0 0 0 vssW
port 39 nsew
flabel metal1 30486 -4531 30686 -4331 0 FreeSans 256 0 0 0 vddW
port 40 nsew
flabel metal1 30380 -5568 30580 -5368 0 FreeSans 256 0 0 0 {la_data_in\[24\]W}
port 28 nsew
flabel metal1 30392 -4922 30592 -4722 0 FreeSans 256 0 0 0 v25W
port 35 nsew
flabel metal1 30392 -6034 30592 -5834 0 FreeSans 256 0 0 0 v18W
port 36 nsew
flabel metal1 32835 -7780 33035 -7580 0 FreeSans 256 0 0 0 {la_data_in\[16\]}
port 18 nsew
flabel metal1 32836 -10180 33036 -9980 0 FreeSans 256 0 0 0 {la_data_in\[17\]}
port 19 nsew
flabel metal1 32836 -12580 33036 -12380 0 FreeSans 256 0 0 0 {la_data_in\[18\]}
port 20 nsew
flabel metal1 32836 -14980 33036 -14780 0 FreeSans 256 0 0 0 {la_data_in\[19\]}
port 21 nsew
flabel metal1 32836 -17380 33036 -17180 0 FreeSans 256 0 0 0 {la_data_in\[20\]}
port 23 nsew
flabel metal1 32836 -19780 33036 -19580 0 FreeSans 256 0 0 0 {la_data_in\[21\]}
port 24 nsew
flabel metal1 32836 -22180 33036 -21980 0 FreeSans 256 0 0 0 {la_data_in\[22\]}
port 25 nsew
flabel metal1 32836 -24580 33036 -24380 0 FreeSans 256 0 0 0 {la_data_in\[23\]}
port 26 nsew
flabel metal1 48596 13343 48796 13543 0 FreeSans 256 0 0 0 {la_data_in\[8\]}
port 0 nsew
flabel metal1 48596 11142 48796 11342 0 FreeSans 256 0 0 0 {la_data_in\[9\]}
port 2 nsew
flabel metal1 48596 8942 48796 9142 0 FreeSans 256 0 0 0 {la_data_in\[10\]}
port 3 nsew
flabel metal1 48596 6742 48796 6942 0 FreeSans 256 0 0 0 {la_data_in\[11\]}
port 8 nsew
flabel metal1 48596 4542 48796 4742 0 FreeSans 256 0 0 0 {la_data_in\[12\]}
port 7 nsew
flabel metal1 48596 2342 48796 2542 0 FreeSans 256 0 0 0 {la_data_in\[13\]}
port 6 nsew
flabel metal1 48575 142 48775 342 0 FreeSans 256 0 0 0 {la_data_in\[14\]}
port 4 nsew
flabel metal1 48596 -2058 48796 -1858 0 FreeSans 256 0 0 0 {la_data_in\[15\]}
port 1 nsew
flabel metal1 48160 -1730 48360 -1530 0 FreeSans 256 0 0 0 {la_data_in\[25\]S}
port 31 nsew
flabel metal1 38140 -24980 38340 -24780 0 FreeSans 256 0 0 0 vssR
port 41 nsew
flabel metal1 45188 -672 45388 -472 0 FreeSans 256 0 0 0 vdd18SI
port 42 nsew
flabel metal1 46052 14708 46252 14908 0 FreeSans 256 0 0 0 vdd25SI
port 43 nsew
flabel metal1 47012 -2526 47212 -2326 0 FreeSans 256 0 0 0 vssSI
port 44 nsew
flabel metal1 58616 62742 58816 62942 0 FreeSans 256 0 0 0 vdd18SO
port 45 nsew
flabel metal1 66980 59150 67180 59350 0 FreeSans 256 0 0 0 vssSO
port 46 nsew
flabel metal1 58950 58735 59150 58935 0 FreeSans 256 0 0 0 Gnd
port 47 nsew
flabel metal1 57552 59058 57752 59258 0 FreeSans 256 0 0 0 vssneg
port 48 nsew
flabel metal1 69890 60551 70090 60751 0 FreeSans 256 0 0 0 {la_data_out\[32\]}
port 50 nsew
flabel metal1 69889 48552 70089 48752 0 FreeSans 256 0 0 0 {la_data_out\[33\]}
port 51 nsew
flabel metal1 69890 36552 70090 36752 0 FreeSans 256 0 0 0 {la_data_out\[34\]}
port 52 nsew
flabel metal1 69890 24552 70090 24752 0 FreeSans 256 0 0 0 {la_data_out\[35\]}
port 53 nsew
flabel metal1 69890 12551 70090 12751 0 FreeSans 256 0 0 0 {la_data_out\[36\]}
port 54 nsew
flabel metal1 69890 552 70090 752 0 FreeSans 256 0 0 0 {la_data_out\[37\]}
port 55 nsew
flabel metal1 69890 -11448 70090 -11248 0 FreeSans 256 0 0 0 {la_data_out\[38\]}
port 56 nsew
flabel metal1 69890 -23448 70090 -23248 0 FreeSans 256 0 0 0 {la_data_out\[39\]}
port 58 nsew
flabel metal2 32180 -1044 32380 -844 0 FreeSans 256 0 0 0 {la_data_in\[25\]B}
port 29 nsew
<< end >>
