magic
tech sky130B
timestamp 1700640568
<< locali >>
rect 2613 1351 2678 3079
rect 2304 1243 2987 1351
rect 2613 -485 2678 1243
<< metal1 >>
rect 2310 -480 2410 -380
rect 2613 -485 2678 1477
<< metal2 >>
rect 2254 1565 2354 1619
rect 2254 1528 2656 1565
rect 2254 1519 2354 1528
rect 2254 -271 2354 -217
rect 2254 -308 2645 -271
rect 2254 -317 2354 -308
<< metal3 >>
rect 2338 3068 2438 3168
rect 2468 3068 2568 3168
rect 2712 3068 2812 3168
rect 2842 3068 2942 3168
rect 2380 1273 2431 3068
rect 2493 1267 2544 3068
rect 2754 1267 2805 3068
rect 2867 1268 2918 3068
use 1T1RLarge  x1
timestamp 1700640568
transform 1 0 2246 0 1 1178
box 8 173 367 1990
use 1T1RLarge  x2
timestamp 1700640568
transform 1 0 2620 0 1 1178
box 8 173 367 1990
use 1T1RLarge  x3
timestamp 1700640568
transform 1 0 2246 0 1 -658
box 8 173 367 1990
use 1T1RLarge  x4
timestamp 1700640568
transform 1 0 2620 0 1 -658
box 8 173 367 1990
<< labels >>
flabel metal1 2310 -480 2410 -380 0 FreeSans 128 0 0 0 VSS
port 6 nsew
flabel metal2 2254 1519 2354 1619 0 FreeSans 128 0 0 0 WL1
port 0 nsew
flabel metal2 2254 -317 2354 -217 0 FreeSans 128 0 0 0 WL2
port 2 nsew
flabel metal3 2712 3068 2812 3168 0 FreeSans 128 0 0 0 SL2
port 5 nsew
flabel metal3 2338 3068 2438 3168 0 FreeSans 128 0 0 0 SL1
port 4 nsew
flabel metal3 2468 3068 2568 3168 0 FreeSans 128 0 0 0 BL1
port 1 nsew
flabel metal3 2842 3068 2942 3168 0 FreeSans 128 0 0 0 BL2
port 3 nsew
<< end >>
