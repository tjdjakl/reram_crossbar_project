magic
tech sky130B
magscale 1 2
timestamp 1700640585
<< metal1 >>
rect -2550 22670 -2350 22870
rect -2644 22278 -2444 22478
rect -2656 21632 -2456 21832
rect -2644 21166 -2444 21366
rect -2552 21006 -2352 21036
rect -2552 20864 -2530 21006
rect -2374 20864 -2352 21006
rect -2552 20836 -2352 20864
rect -74 20488 -64 20630
rect 76 20488 86 20630
rect -200 19420 0 19620
rect 1440 19416 1640 19616
rect 870 18666 880 18786
rect 1040 18666 1050 18786
rect -80 18106 -70 18214
rect 82 18106 92 18214
rect -200 17020 0 17220
rect 1440 17016 1640 17216
rect 868 16258 878 16378
rect 1038 16258 1048 16378
rect -80 15702 -70 15810
rect 82 15702 92 15810
rect -200 14620 0 14820
rect 1440 14616 1640 14816
rect 870 13868 880 13988
rect 1040 13868 1050 13988
rect -78 13296 -68 13404
rect 84 13296 94 13404
rect -200 12220 0 12420
rect 1440 12216 1640 12416
rect 866 11464 876 11584
rect 1036 11464 1046 11584
rect -80 10884 -70 10992
rect 82 10884 92 10992
rect -200 9820 0 10020
rect 1440 9816 1640 10016
rect 872 9066 882 9186
rect 1042 9066 1052 9186
rect -78 8498 -68 8606
rect 84 8498 94 8606
rect -200 7420 0 7620
rect 1440 7416 1640 7616
rect 866 6666 876 6786
rect 1036 6666 1046 6786
rect -84 6092 -74 6200
rect 78 6092 88 6200
rect -200 5020 0 5220
rect 1440 5016 1640 5216
rect 858 4264 868 4384
rect 1028 4264 1038 4384
rect -80 3720 -70 3828
rect 82 3720 92 3828
rect -200 2620 0 2820
rect 1440 2616 1640 2816
rect 868 1868 878 1988
rect 1038 1868 1048 1988
<< via1 >>
rect -2530 20864 -2374 21006
rect -64 20488 76 20630
rect 880 18666 1040 18786
rect -70 18106 82 18214
rect 878 16258 1038 16378
rect -70 15702 82 15810
rect 880 13868 1040 13988
rect -68 13296 84 13404
rect 876 11464 1036 11584
rect -70 10884 82 10992
rect 882 9066 1042 9186
rect -68 8498 84 8606
rect 876 6666 1036 6786
rect -74 6092 78 6200
rect 868 4264 1028 4384
rect -70 3720 82 3828
rect 878 1868 1038 1988
<< metal2 >>
rect -2530 21006 -2374 21016
rect -2530 20854 -2374 20864
rect -64 20630 76 21770
rect -64 18224 76 20488
rect 880 20972 1038 20988
rect 880 20860 886 20972
rect 1036 20860 1038 20972
rect 880 18796 1038 20860
rect 880 18786 1040 18796
rect 878 18666 880 18736
rect 878 18656 1040 18666
rect -70 18214 82 18224
rect -70 18096 82 18106
rect -64 15820 76 18096
rect 878 16378 1038 18656
rect -70 15810 82 15820
rect -70 15692 82 15702
rect -64 13414 76 15692
rect 878 13998 1038 16258
rect 878 13988 1040 13998
rect 878 13868 880 13988
rect 878 13858 1040 13868
rect -68 13404 84 13414
rect -68 13286 84 13296
rect -64 11002 76 13286
rect 878 11594 1038 13858
rect 876 11584 1038 11594
rect 1036 11464 1038 11584
rect 876 11454 1038 11464
rect -70 10992 82 11002
rect -70 10874 82 10884
rect -64 8616 76 10874
rect 878 9196 1038 11454
rect 878 9186 1042 9196
rect 878 9066 882 9186
rect 878 9056 1042 9066
rect -68 8606 84 8616
rect -68 8488 84 8498
rect -64 6210 76 8488
rect 878 6796 1038 9056
rect 876 6786 1038 6796
rect 1036 6666 1038 6786
rect 876 6656 1038 6666
rect -74 6200 78 6210
rect -74 6082 78 6092
rect -64 3838 76 6082
rect 878 4394 1038 6656
rect 868 4384 1038 4394
rect 1028 4264 1038 4384
rect 868 4254 1038 4264
rect -70 3828 82 3838
rect -70 3710 82 3720
rect 878 1988 1038 4254
rect 878 1858 1038 1868
<< via2 >>
rect -2530 20864 -2374 21006
rect 886 20860 1036 20972
<< metal3 >>
rect -2540 21006 -2364 21011
rect -2540 20864 -2530 21006
rect -2374 21004 -2364 21006
rect -2374 20977 1036 21004
rect -2374 20972 1046 20977
rect -2374 20864 886 20972
rect -2540 20859 -2364 20864
rect 876 20860 886 20864
rect 1036 20860 1046 20972
rect 876 20855 1046 20860
use Buffer  x1
timestamp 1700618825
transform 1 0 -2058 0 1 17240
box 1858 1360 3698 3442
use Buffer  x2
timestamp 1700618825
transform 1 0 -2058 0 1 14840
box 1858 1360 3698 3442
use Buffer  x3
timestamp 1700618825
transform 1 0 -2058 0 1 12440
box 1858 1360 3698 3442
use Buffer  x4
timestamp 1700618825
transform 1 0 -2058 0 1 10040
box 1858 1360 3698 3442
use Buffer  x5
timestamp 1700618825
transform 1 0 -2058 0 1 7640
box 1858 1360 3698 3442
use Buffer  x6
timestamp 1700618825
transform 1 0 -2058 0 1 5240
box 1858 1360 3698 3442
use Buffer  x7
timestamp 1700618825
transform 1 0 -2058 0 1 2840
box 1858 1360 3698 3442
use Buffer  x8
timestamp 1700618825
transform 1 0 -2058 0 1 440
box 1858 1360 3698 3442
use 2-1MUX  x9
timestamp 1700640585
transform 1 0 -1720 0 1 20180
box -936 600 1824 2716
<< labels >>
flabel metal1 -2550 22670 -2350 22870 0 FreeSans 256 0 0 0 VDD
port 17 nsew
flabel metal1 -2552 20836 -2352 21036 0 FreeSans 256 0 0 0 VSS
port 18 nsew
flabel metal1 -200 19420 0 19620 0 FreeSans 256 0 0 0 WL_LA_IN1
port 0 nsew
flabel metal1 -200 17020 0 17220 0 FreeSans 256 0 0 0 WL_LA_IN2
port 1 nsew
flabel metal1 -200 14620 0 14820 0 FreeSans 256 0 0 0 WL_LA_IN3
port 2 nsew
flabel metal1 -200 12220 0 12420 0 FreeSans 256 0 0 0 WL_LA_IN4
port 3 nsew
flabel metal1 -200 9820 0 10020 0 FreeSans 256 0 0 0 WL_LA_IN5
port 4 nsew
flabel metal1 -200 7420 0 7620 0 FreeSans 256 0 0 0 WL_LA_IN6
port 5 nsew
flabel metal1 -200 5020 0 5220 0 FreeSans 256 0 0 0 WL_LA_IN7
port 6 nsew
flabel metal1 -200 2620 0 2820 0 FreeSans 256 0 0 0 WL_LA_IN8
port 8 nsew
flabel metal1 1440 19416 1640 19616 0 FreeSans 256 0 0 0 WL_IN1
port 9 nsew
flabel metal1 1440 17016 1640 17216 0 FreeSans 256 0 0 0 WL_IN2
port 10 nsew
flabel metal1 1440 14616 1640 14816 0 FreeSans 256 0 0 0 WL_IN3
port 11 nsew
flabel metal1 1440 12216 1640 12416 0 FreeSans 256 0 0 0 WL_IN4
port 12 nsew
flabel metal1 1440 9816 1640 10016 0 FreeSans 256 0 0 0 WL_IN5
port 13 nsew
flabel metal1 1440 7416 1640 7616 0 FreeSans 256 0 0 0 WL_IN6
port 14 nsew
flabel metal1 1440 5016 1640 5216 0 FreeSans 256 0 0 0 WL_IN7
port 15 nsew
flabel metal1 1440 2616 1640 2816 0 FreeSans 256 0 0 0 WL_IN8
port 16 nsew
flabel metal1 -2656 21632 -2456 21832 0 FreeSans 256 0 0 0 Write_Select
port 19 nsew
flabel metal1 -2644 22278 -2444 22478 0 FreeSans 256 0 0 0 Write_Voltage
port 20 nsew
flabel metal1 -2644 21166 -2444 21366 0 FreeSans 256 0 0 0 Form_Voltage
port 22 nsew
<< end >>
