magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect -38 261 2614 582
<< pwell >>
rect 1408 157 1769 201
rect 2298 157 2575 203
rect 1 21 2575 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 151 47 181 131
rect 235 47 265 131
rect 319 47 349 131
rect 513 47 543 131
rect 701 47 731 131
rect 785 47 815 131
rect 973 47 1003 131
rect 1057 47 1087 131
rect 1129 47 1159 131
rect 1317 47 1347 131
rect 1389 47 1419 131
rect 1484 47 1514 175
rect 1663 47 1693 175
rect 1785 47 1815 131
rect 1857 47 1887 131
rect 1953 47 1983 131
rect 2067 47 2097 131
rect 2279 47 2309 131
rect 2374 47 2404 177
rect 2467 47 2497 177
<< scpmoshvt >>
rect 79 369 109 497
rect 163 369 193 497
rect 235 369 265 497
rect 319 369 349 497
rect 507 369 537 497
rect 695 369 725 497
rect 779 369 809 497
rect 967 413 997 497
rect 1051 413 1081 497
rect 1153 413 1183 497
rect 1281 413 1311 497
rect 1379 413 1409 497
rect 1495 329 1525 497
rect 1567 329 1597 497
rect 1693 413 1723 497
rect 1781 413 1811 497
rect 1903 413 1933 497
rect 2091 413 2121 497
rect 2279 360 2309 488
rect 2374 297 2404 497
rect 2467 297 2497 497
<< ndiff >>
rect 1434 131 1484 175
rect 27 103 79 131
rect 27 69 35 103
rect 69 69 79 103
rect 27 47 79 69
rect 109 47 151 131
rect 181 93 235 131
rect 181 59 191 93
rect 225 59 235 93
rect 181 47 235 59
rect 265 47 319 131
rect 349 93 407 131
rect 349 59 365 93
rect 399 59 407 93
rect 349 47 407 59
rect 461 105 513 131
rect 461 71 469 105
rect 503 71 513 105
rect 461 47 513 71
rect 543 93 595 131
rect 543 59 553 93
rect 587 59 595 93
rect 543 47 595 59
rect 649 105 701 131
rect 649 71 657 105
rect 691 71 701 105
rect 649 47 701 71
rect 731 89 785 131
rect 731 55 741 89
rect 775 55 785 89
rect 731 47 785 55
rect 815 101 867 131
rect 815 67 825 101
rect 859 67 867 101
rect 815 47 867 67
rect 921 101 973 131
rect 921 67 929 101
rect 963 67 973 101
rect 921 47 973 67
rect 1003 101 1057 131
rect 1003 67 1013 101
rect 1047 67 1057 101
rect 1003 47 1057 67
rect 1087 47 1129 131
rect 1159 93 1211 131
rect 1159 59 1169 93
rect 1203 59 1211 93
rect 1159 47 1211 59
rect 1265 119 1317 131
rect 1265 85 1273 119
rect 1307 85 1317 119
rect 1265 47 1317 85
rect 1347 47 1389 131
rect 1419 89 1484 131
rect 1419 55 1431 89
rect 1465 55 1484 89
rect 1419 47 1484 55
rect 1514 47 1663 175
rect 1693 131 1743 175
rect 2324 131 2374 177
rect 1693 89 1785 131
rect 1693 55 1709 89
rect 1743 55 1785 89
rect 1693 47 1785 55
rect 1815 47 1857 131
rect 1887 47 1953 131
rect 1983 89 2067 131
rect 1983 55 2023 89
rect 2057 55 2067 89
rect 1983 47 2067 55
rect 2097 101 2173 131
rect 2097 67 2131 101
rect 2165 67 2173 101
rect 2097 47 2173 67
rect 2227 102 2279 131
rect 2227 68 2235 102
rect 2269 68 2279 102
rect 2227 47 2279 68
rect 2309 89 2374 131
rect 2309 55 2330 89
rect 2364 55 2374 89
rect 2309 47 2374 55
rect 2404 157 2467 177
rect 2404 123 2423 157
rect 2457 123 2467 157
rect 2404 89 2467 123
rect 2404 55 2423 89
rect 2457 55 2467 89
rect 2404 47 2467 55
rect 2497 161 2549 177
rect 2497 127 2507 161
rect 2541 127 2549 161
rect 2497 93 2549 127
rect 2497 59 2507 93
rect 2541 59 2549 93
rect 2497 47 2549 59
<< pdiff >>
rect 27 431 79 497
rect 27 397 35 431
rect 69 397 79 431
rect 27 369 79 397
rect 109 489 163 497
rect 109 455 119 489
rect 153 455 163 489
rect 109 369 163 455
rect 193 369 235 497
rect 265 411 319 497
rect 265 377 275 411
rect 309 377 319 411
rect 265 369 319 377
rect 349 485 401 497
rect 349 451 359 485
rect 393 451 401 485
rect 349 369 401 451
rect 455 415 507 497
rect 455 381 463 415
rect 497 381 507 415
rect 455 369 507 381
rect 537 485 589 497
rect 537 451 547 485
rect 581 451 589 485
rect 537 369 589 451
rect 643 449 695 497
rect 643 415 651 449
rect 685 415 695 449
rect 643 369 695 415
rect 725 489 779 497
rect 725 455 735 489
rect 769 455 779 489
rect 725 369 779 455
rect 809 477 861 497
rect 809 443 819 477
rect 853 443 861 477
rect 809 369 861 443
rect 915 477 967 497
rect 915 443 923 477
rect 957 443 967 477
rect 915 413 967 443
rect 997 477 1051 497
rect 997 443 1007 477
rect 1041 443 1051 477
rect 997 413 1051 443
rect 1081 413 1153 497
rect 1183 489 1281 497
rect 1183 455 1205 489
rect 1239 455 1281 489
rect 1183 413 1281 455
rect 1311 474 1379 497
rect 1311 440 1326 474
rect 1360 440 1379 474
rect 1311 413 1379 440
rect 1409 489 1495 497
rect 1409 455 1428 489
rect 1462 455 1495 489
rect 1409 413 1495 455
rect 1445 329 1495 413
rect 1525 329 1567 497
rect 1597 475 1693 497
rect 1597 441 1637 475
rect 1671 441 1693 475
rect 1597 413 1693 441
rect 1723 413 1781 497
rect 1811 489 1903 497
rect 1811 455 1848 489
rect 1882 455 1903 489
rect 1811 413 1903 455
rect 1933 474 1985 497
rect 1933 440 1943 474
rect 1977 440 1985 474
rect 1933 413 1985 440
rect 2039 485 2091 497
rect 2039 451 2047 485
rect 2081 451 2091 485
rect 2039 413 2091 451
rect 2121 474 2173 497
rect 2324 488 2374 497
rect 2121 440 2131 474
rect 2165 440 2173 474
rect 2121 413 2173 440
rect 2227 476 2279 488
rect 2227 442 2235 476
rect 2269 442 2279 476
rect 1597 329 1647 413
rect 2227 408 2279 442
rect 2227 374 2235 408
rect 2269 374 2279 408
rect 2227 360 2279 374
rect 2309 476 2374 488
rect 2309 442 2330 476
rect 2364 442 2374 476
rect 2309 408 2374 442
rect 2309 374 2330 408
rect 2364 374 2374 408
rect 2309 360 2374 374
rect 2324 297 2374 360
rect 2404 485 2467 497
rect 2404 451 2423 485
rect 2457 451 2467 485
rect 2404 417 2467 451
rect 2404 383 2423 417
rect 2457 383 2467 417
rect 2404 349 2467 383
rect 2404 315 2423 349
rect 2457 315 2467 349
rect 2404 297 2467 315
rect 2497 485 2549 497
rect 2497 451 2507 485
rect 2541 451 2549 485
rect 2497 417 2549 451
rect 2497 383 2507 417
rect 2541 383 2549 417
rect 2497 349 2549 383
rect 2497 315 2507 349
rect 2541 315 2549 349
rect 2497 297 2549 315
<< ndiffc >>
rect 35 69 69 103
rect 191 59 225 93
rect 365 59 399 93
rect 469 71 503 105
rect 553 59 587 93
rect 657 71 691 105
rect 741 55 775 89
rect 825 67 859 101
rect 929 67 963 101
rect 1013 67 1047 101
rect 1169 59 1203 93
rect 1273 85 1307 119
rect 1431 55 1465 89
rect 1709 55 1743 89
rect 2023 55 2057 89
rect 2131 67 2165 101
rect 2235 68 2269 102
rect 2330 55 2364 89
rect 2423 123 2457 157
rect 2423 55 2457 89
rect 2507 127 2541 161
rect 2507 59 2541 93
<< pdiffc >>
rect 35 397 69 431
rect 119 455 153 489
rect 275 377 309 411
rect 359 451 393 485
rect 463 381 497 415
rect 547 451 581 485
rect 651 415 685 449
rect 735 455 769 489
rect 819 443 853 477
rect 923 443 957 477
rect 1007 443 1041 477
rect 1205 455 1239 489
rect 1326 440 1360 474
rect 1428 455 1462 489
rect 1637 441 1671 475
rect 1848 455 1882 489
rect 1943 440 1977 474
rect 2047 451 2081 485
rect 2131 440 2165 474
rect 2235 442 2269 476
rect 2235 374 2269 408
rect 2330 442 2364 476
rect 2330 374 2364 408
rect 2423 451 2457 485
rect 2423 383 2457 417
rect 2423 315 2457 349
rect 2507 451 2541 485
rect 2507 383 2541 417
rect 2507 315 2541 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 235 497 265 523
rect 319 497 349 523
rect 507 497 537 523
rect 695 497 725 523
rect 779 497 809 523
rect 967 497 997 523
rect 1051 497 1081 523
rect 1153 497 1183 523
rect 1281 497 1311 523
rect 1379 497 1409 523
rect 1495 497 1525 523
rect 1567 497 1597 523
rect 1693 497 1723 523
rect 1781 497 1811 523
rect 1903 497 1933 523
rect 2091 497 2121 523
rect 967 398 997 413
rect 79 354 109 369
rect 48 324 109 354
rect 48 265 78 324
rect 163 283 193 369
rect 21 249 78 265
rect 21 215 34 249
rect 68 215 78 249
rect 120 267 193 283
rect 120 233 130 267
rect 164 253 193 267
rect 164 233 181 253
rect 120 217 181 233
rect 235 219 265 369
rect 319 265 349 369
rect 507 265 537 369
rect 695 354 725 369
rect 683 324 725 354
rect 683 284 713 324
rect 779 284 809 369
rect 908 368 997 398
rect 1051 381 1081 413
rect 1153 381 1183 413
rect 908 284 938 368
rect 1039 365 1093 381
rect 1039 331 1049 365
rect 1083 331 1093 365
rect 1039 315 1093 331
rect 1153 365 1229 381
rect 1153 331 1185 365
rect 1219 331 1229 365
rect 1153 315 1229 331
rect 659 268 713 284
rect 319 249 438 265
rect 21 199 78 215
rect 48 176 78 199
rect 48 146 109 176
rect 79 131 109 146
rect 151 131 181 217
rect 223 203 277 219
rect 223 169 233 203
rect 267 169 277 203
rect 223 153 277 169
rect 319 215 373 249
rect 407 215 438 249
rect 319 199 438 215
rect 480 249 543 265
rect 480 215 490 249
rect 524 215 543 249
rect 659 234 669 268
rect 703 234 713 268
rect 659 218 713 234
rect 755 268 812 284
rect 755 234 765 268
rect 799 234 812 268
rect 755 218 812 234
rect 854 268 938 284
rect 854 234 864 268
rect 898 248 938 268
rect 898 234 1087 248
rect 854 218 1087 234
rect 480 199 543 215
rect 235 131 265 153
rect 319 131 349 199
rect 513 131 543 199
rect 683 176 713 218
rect 782 176 812 218
rect 683 146 731 176
rect 782 146 1003 176
rect 701 131 731 146
rect 785 131 815 146
rect 973 131 1003 146
rect 1057 131 1087 218
rect 1153 213 1183 315
rect 1281 273 1311 413
rect 1379 369 1409 413
rect 1353 353 1409 369
rect 1353 319 1363 353
rect 1397 319 1409 353
rect 2279 488 2309 523
rect 2374 497 2404 523
rect 2467 497 2497 523
rect 1693 381 1723 413
rect 1685 365 1739 381
rect 1685 345 1695 365
rect 1663 331 1695 345
rect 1729 331 1739 365
rect 1353 303 1409 319
rect 1245 263 1311 273
rect 1245 229 1261 263
rect 1295 229 1311 263
rect 1379 273 1409 303
rect 1379 243 1419 273
rect 1495 265 1525 329
rect 1245 219 1311 229
rect 1129 203 1195 213
rect 1129 169 1145 203
rect 1179 169 1195 203
rect 1129 159 1195 169
rect 1281 176 1311 219
rect 1129 131 1159 159
rect 1281 146 1347 176
rect 1317 131 1347 146
rect 1389 131 1419 243
rect 1461 249 1525 265
rect 1461 215 1471 249
rect 1505 215 1525 249
rect 1461 199 1525 215
rect 1567 265 1597 329
rect 1663 315 1739 331
rect 1781 325 1811 413
rect 1903 397 1933 413
rect 1903 367 1983 397
rect 1929 343 1983 367
rect 2091 365 2121 413
rect 1567 249 1621 265
rect 1567 215 1577 249
rect 1611 215 1621 249
rect 1567 199 1621 215
rect 1484 175 1514 199
rect 1663 175 1693 315
rect 1781 295 1887 325
rect 1761 235 1815 251
rect 1761 201 1771 235
rect 1805 201 1815 235
rect 1761 185 1815 201
rect 1785 131 1815 185
rect 1857 237 1887 295
rect 1929 309 1939 343
rect 1973 309 1983 343
rect 2031 355 2121 365
rect 2031 321 2047 355
rect 2081 341 2121 355
rect 2279 341 2309 360
rect 2081 321 2309 341
rect 2031 311 2309 321
rect 1929 293 1983 309
rect 1857 221 1911 237
rect 1857 187 1867 221
rect 1901 187 1911 221
rect 1857 171 1911 187
rect 1857 131 1887 171
rect 1953 131 1983 293
rect 2043 203 2097 311
rect 2043 169 2053 203
rect 2087 169 2097 203
rect 2043 153 2097 169
rect 2067 131 2097 153
rect 2279 131 2309 311
rect 2374 265 2404 297
rect 2467 265 2497 297
rect 2351 249 2497 265
rect 2351 215 2361 249
rect 2395 215 2497 249
rect 2351 199 2497 215
rect 2374 177 2404 199
rect 2467 177 2497 199
rect 79 21 109 47
rect 151 21 181 47
rect 235 21 265 47
rect 319 21 349 47
rect 513 21 543 47
rect 701 21 731 47
rect 785 21 815 47
rect 973 21 1003 47
rect 1057 21 1087 47
rect 1129 21 1159 47
rect 1317 21 1347 47
rect 1389 21 1419 47
rect 1484 21 1514 47
rect 1663 21 1693 47
rect 1785 21 1815 47
rect 1857 21 1887 47
rect 1953 21 1983 47
rect 2067 21 2097 47
rect 2279 21 2309 47
rect 2374 21 2404 47
rect 2467 21 2497 47
<< polycont >>
rect 34 215 68 249
rect 130 233 164 267
rect 1049 331 1083 365
rect 1185 331 1219 365
rect 233 169 267 203
rect 373 215 407 249
rect 490 215 524 249
rect 669 234 703 268
rect 765 234 799 268
rect 864 234 898 268
rect 1363 319 1397 353
rect 1695 331 1729 365
rect 1261 229 1295 263
rect 1145 169 1179 203
rect 1471 215 1505 249
rect 1577 215 1611 249
rect 1771 201 1805 235
rect 1939 309 1973 343
rect 2047 321 2081 355
rect 1867 187 1901 221
rect 2053 169 2087 203
rect 2361 215 2395 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 17 431 69 493
rect 103 489 157 527
rect 103 455 119 489
rect 153 455 157 489
rect 103 439 157 455
rect 191 485 409 493
rect 191 451 359 485
rect 393 451 409 485
rect 17 397 35 431
rect 191 405 225 451
rect 454 417 504 493
rect 538 485 597 527
rect 538 451 547 485
rect 581 451 597 485
rect 719 489 785 527
rect 538 428 597 451
rect 651 449 685 465
rect 719 455 735 489
rect 769 455 785 489
rect 819 477 888 493
rect 69 397 225 405
rect 17 369 225 397
rect 259 411 339 417
rect 259 377 275 411
rect 309 377 339 411
rect 259 369 339 377
rect 17 249 68 335
rect 17 215 34 249
rect 17 153 68 215
rect 108 267 164 335
rect 108 255 130 267
rect 108 221 121 255
rect 155 221 164 233
rect 108 153 164 221
rect 210 203 267 335
rect 210 169 233 203
rect 210 153 267 169
rect 301 323 339 369
rect 301 289 305 323
rect 301 142 339 289
rect 373 415 504 417
rect 373 381 463 415
rect 497 381 504 415
rect 853 443 888 477
rect 819 427 888 443
rect 651 400 685 415
rect 651 398 797 400
rect 373 354 504 381
rect 373 249 440 354
rect 581 323 617 392
rect 651 391 799 398
rect 651 366 765 391
rect 747 357 765 366
rect 407 215 440 249
rect 474 255 540 320
rect 474 221 489 255
rect 523 249 540 255
rect 474 215 490 221
rect 524 215 540 249
rect 581 268 713 323
rect 581 234 669 268
rect 703 234 713 268
rect 373 181 440 215
rect 581 211 713 234
rect 747 268 799 357
rect 747 234 765 268
rect 373 143 504 181
rect 581 145 620 211
rect 747 177 799 234
rect 301 141 335 142
rect 299 133 335 141
rect 295 132 335 133
rect 295 129 334 132
rect 292 127 333 129
rect 289 126 333 127
rect 288 124 333 126
rect 286 123 332 124
rect 284 122 332 123
rect 281 121 332 122
rect 279 120 332 121
rect 276 119 332 120
rect 17 103 140 119
rect 17 69 35 103
rect 69 69 140 103
rect 17 17 140 69
rect 174 115 330 119
rect 174 111 328 115
rect 174 93 325 111
rect 174 59 191 93
rect 225 59 325 93
rect 174 51 325 59
rect 365 93 418 109
rect 399 59 418 93
rect 365 17 418 59
rect 452 105 504 143
rect 654 143 799 177
rect 833 284 888 427
rect 923 477 966 493
rect 957 443 966 477
rect 923 323 966 443
rect 1007 477 1151 493
rect 1041 443 1151 477
rect 1189 489 1266 527
rect 1189 455 1205 489
rect 1239 455 1266 489
rect 1321 474 1364 490
rect 1007 427 1151 443
rect 1075 365 1083 391
rect 1041 331 1049 357
rect 923 318 949 323
rect 932 289 949 318
rect 1041 315 1083 331
rect 833 268 898 284
rect 833 255 864 268
rect 833 221 857 255
rect 891 221 898 234
rect 833 218 898 221
rect 452 71 469 105
rect 503 71 504 105
rect 452 51 504 71
rect 538 93 620 111
rect 538 59 553 93
rect 587 59 620 93
rect 538 17 620 59
rect 654 105 691 143
rect 833 117 867 218
rect 932 184 966 289
rect 1117 279 1151 427
rect 1321 440 1326 474
rect 1360 440 1364 474
rect 1321 421 1364 440
rect 1412 489 1603 527
rect 1412 455 1428 489
rect 1462 455 1603 489
rect 1412 425 1603 455
rect 1637 475 1798 492
rect 1671 441 1798 475
rect 1832 489 1898 527
rect 1832 455 1848 489
rect 1882 455 1898 489
rect 1832 447 1898 455
rect 1932 474 1993 490
rect 1637 425 1798 441
rect 1185 387 1364 421
rect 1764 413 1798 425
rect 1932 440 1943 474
rect 1977 440 1993 474
rect 2031 485 2097 527
rect 2031 451 2047 485
rect 2081 451 2097 485
rect 2031 447 2097 451
rect 2131 474 2183 493
rect 1932 413 1993 440
rect 2165 440 2183 474
rect 1185 365 1219 387
rect 1447 357 1512 391
rect 1546 357 1627 391
rect 1185 315 1219 331
rect 1328 323 1363 353
rect 1362 319 1363 323
rect 1397 319 1413 353
rect 1447 334 1627 357
rect 1362 289 1413 319
rect 1017 263 1295 279
rect 1017 255 1261 263
rect 654 71 657 105
rect 654 51 691 71
rect 725 89 791 109
rect 725 55 741 89
rect 775 55 791 89
rect 725 17 791 55
rect 825 101 867 117
rect 859 67 867 101
rect 825 51 867 67
rect 901 101 966 184
rect 901 67 929 101
rect 963 67 966 101
rect 901 51 966 67
rect 1000 245 1261 255
rect 1000 101 1088 245
rect 1471 255 1543 265
rect 1295 249 1543 255
rect 1295 229 1471 249
rect 1261 215 1471 229
rect 1505 215 1543 249
rect 1129 169 1145 203
rect 1179 169 1195 203
rect 1261 195 1543 215
rect 1577 249 1627 334
rect 1611 215 1627 249
rect 1685 365 1730 381
rect 1764 379 2097 413
rect 1685 331 1695 365
rect 1729 331 1730 365
rect 2031 355 2097 379
rect 1685 255 1730 331
rect 1776 343 1989 345
rect 1776 323 1939 343
rect 1776 289 1788 323
rect 1822 309 1939 323
rect 1973 309 1989 343
rect 2031 321 2047 355
rect 2081 321 2097 355
rect 1822 289 1827 309
rect 1776 285 1827 289
rect 2131 273 2183 440
rect 1685 221 1696 255
rect 1685 215 1730 221
rect 1764 235 1821 251
rect 1129 161 1195 169
rect 1577 181 1627 215
rect 1764 201 1771 235
rect 1805 201 1821 235
rect 1764 181 1821 201
rect 1129 127 1307 161
rect 1000 67 1013 101
rect 1047 67 1088 101
rect 1257 119 1307 127
rect 1000 51 1088 67
rect 1122 59 1169 93
rect 1203 59 1219 93
rect 1122 17 1219 59
rect 1257 85 1273 119
rect 1257 51 1307 85
rect 1341 89 1543 161
rect 1577 144 1821 181
rect 1864 239 2183 273
rect 1864 221 1906 239
rect 1864 187 1867 221
rect 1901 187 1906 221
rect 1864 171 1906 187
rect 1942 169 2053 203
rect 2087 169 2103 203
rect 1942 157 2103 169
rect 1942 109 1982 157
rect 2137 117 2183 239
rect 1341 55 1431 89
rect 1465 55 1543 89
rect 1693 89 1982 109
rect 1693 55 1709 89
rect 1743 55 1982 89
rect 2023 89 2073 109
rect 2057 55 2073 89
rect 1341 17 1543 55
rect 2023 17 2073 55
rect 2115 101 2183 117
rect 2115 67 2131 101
rect 2165 67 2183 101
rect 2115 51 2183 67
rect 2217 476 2269 493
rect 2217 442 2235 476
rect 2217 408 2269 442
rect 2217 374 2235 408
rect 2217 265 2269 374
rect 2314 476 2364 527
rect 2314 442 2330 476
rect 2314 408 2364 442
rect 2314 374 2330 408
rect 2314 358 2364 374
rect 2407 485 2473 490
rect 2407 451 2423 485
rect 2457 451 2473 485
rect 2407 417 2473 451
rect 2407 383 2423 417
rect 2457 383 2473 417
rect 2407 349 2473 383
rect 2407 315 2423 349
rect 2457 315 2473 349
rect 2407 299 2473 315
rect 2507 485 2559 527
rect 2541 451 2559 485
rect 2507 417 2559 451
rect 2541 383 2559 417
rect 2507 349 2559 383
rect 2541 315 2559 349
rect 2507 299 2559 315
rect 2217 249 2395 265
rect 2217 215 2361 249
rect 2217 199 2395 215
rect 2217 102 2269 199
rect 2429 165 2473 299
rect 2217 68 2235 102
rect 2217 51 2269 68
rect 2314 89 2373 165
rect 2314 55 2330 89
rect 2364 55 2373 89
rect 2314 17 2373 55
rect 2407 157 2473 165
rect 2407 123 2423 157
rect 2457 123 2473 157
rect 2407 89 2473 123
rect 2407 55 2423 89
rect 2457 55 2473 89
rect 2407 51 2473 55
rect 2507 161 2559 177
rect 2541 127 2559 161
rect 2507 93 2559 127
rect 2541 59 2559 93
rect 2507 17 2559 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 121 233 130 255
rect 130 233 155 255
rect 121 221 155 233
rect 305 289 339 323
rect 765 357 799 391
rect 489 249 523 255
rect 489 221 490 249
rect 490 221 523 249
rect 1041 365 1075 391
rect 1041 357 1049 365
rect 1049 357 1075 365
rect 949 289 983 323
rect 857 234 864 255
rect 864 234 891 255
rect 857 221 891 234
rect 1512 357 1546 391
rect 1328 289 1362 323
rect 1788 289 1822 323
rect 1696 221 1730 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
<< metal1 >>
rect 0 561 2576 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 0 496 2576 527
rect 753 391 811 397
rect 753 357 765 391
rect 799 388 811 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 799 360 1041 388
rect 799 357 811 360
rect 753 351 811 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1500 391 1558 397
rect 1500 388 1512 391
rect 1075 360 1512 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1500 357 1512 360
rect 1546 357 1558 391
rect 1500 351 1558 357
rect 293 323 351 329
rect 293 289 305 323
rect 339 320 351 323
rect 937 323 995 329
rect 937 320 949 323
rect 339 292 949 320
rect 339 289 351 292
rect 293 283 351 289
rect 937 289 949 292
rect 983 289 995 323
rect 937 283 995 289
rect 1316 323 1374 329
rect 1316 289 1328 323
rect 1362 320 1374 323
rect 1776 323 1834 329
rect 1776 320 1788 323
rect 1362 292 1788 320
rect 1362 289 1374 292
rect 1316 283 1374 289
rect 1776 289 1788 292
rect 1822 289 1834 323
rect 1776 283 1834 289
rect 109 255 167 261
rect 109 221 121 255
rect 155 252 167 255
rect 477 255 535 261
rect 477 252 489 255
rect 155 224 489 252
rect 155 221 167 224
rect 109 215 167 221
rect 477 221 489 224
rect 523 221 535 255
rect 477 215 535 221
rect 845 255 903 261
rect 845 221 857 255
rect 891 252 903 255
rect 1684 255 1742 261
rect 1684 252 1696 255
rect 891 224 1696 252
rect 891 221 903 224
rect 845 215 903 221
rect 1684 221 1696 224
rect 1730 221 1742 255
rect 1684 215 1742 221
rect 0 17 2576 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
rect 0 -48 2576 -17
<< labels >>
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 SCD
port 3 nsew signal input
flabel locali s 581 357 615 391 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 213 289 247 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 SCD
port 3 nsew signal input
flabel locali s 1328 289 1362 323 0 FreeSans 200 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 SCE
port 4 nsew signal input
flabel locali s 213 153 247 187 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 581 153 615 187 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2439 357 2473 391 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2439 425 2473 459 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2439 221 2473 255 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2439 153 2473 187 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2439 85 2473 119 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2439 289 2473 323 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 sdfstp_2
flabel comment s 1168 291 1168 291 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 2069 226 2069 226 0 FreeSans 200 0 0 0 no_jumper_check
rlabel locali s 474 215 540 320 1 SCE
port 4 nsew signal input
rlabel metal1 s 477 252 535 261 1 SCE
port 4 nsew signal input
rlabel metal1 s 477 215 535 224 1 SCE
port 4 nsew signal input
rlabel metal1 s 109 252 167 261 1 SCE
port 4 nsew signal input
rlabel metal1 s 109 224 535 252 1 SCE
port 4 nsew signal input
rlabel metal1 s 109 215 167 224 1 SCE
port 4 nsew signal input
rlabel locali s 1776 309 1989 345 1 SET_B
port 5 nsew signal input
rlabel locali s 1776 285 1827 309 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1776 320 1834 329 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1776 283 1834 292 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 320 1374 329 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 292 1834 320 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 283 1374 292 1 SET_B
port 5 nsew signal input
rlabel metal1 s 0 -48 2576 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2576 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2576 544
string GDS_END 304536
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 284032
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 12.880 2.720 
<< end >>
