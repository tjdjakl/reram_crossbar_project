magic
tech sky130B
timestamp 1700618825
<< locali >>
rect 1031 3888 1094 4797
rect 1378 3751 1441 4797
rect 1727 3888 1788 4797
rect 745 3641 2074 3751
rect 1034 2595 1095 2723
rect 1378 2595 1441 3641
rect 745 2501 2074 2595
rect 1014 1592 1095 2501
rect 1034 1456 1095 1592
rect 1378 1456 1441 2501
rect 1727 1593 1788 2501
rect 745 1346 2074 1456
rect 1378 300 1441 1346
<< metal1 >>
rect 1371 3751 1444 3888
rect 1034 1433 1095 2737
rect 1383 2732 1444 3751
rect 1372 2595 1444 2732
rect 1383 1593 1444 2595
rect 1731 1593 1792 2598
rect 1374 1456 1444 1593
rect 1383 437 1444 1456
rect 759 310 859 410
rect 1378 300 1445 437
<< metal2 >>
rect 689 3935 789 4035
rect 1019 3949 1440 4021
rect 689 2779 789 2879
rect 1016 2794 1437 2866
rect 689 1640 789 1740
rect 1011 1654 1432 1726
rect 689 484 789 584
rect 980 499 1401 571
<< metal3 >>
rect 778 4780 878 4880
rect 911 4780 1011 4880
rect 1125 4780 1225 4880
rect 1258 4780 1358 4880
rect 1474 4780 1574 4880
rect 1607 4780 1707 4880
rect 1821 4780 1921 4880
rect 1954 4780 2054 4880
rect 787 2520 866 3737
rect 919 1393 998 4780
rect 1134 2521 1213 3738
rect 1266 1382 1345 4780
rect 1483 2523 1562 3740
rect 1615 1381 1694 4780
rect 1830 2527 1909 3744
rect 1962 1388 2041 4780
use 4T4R  x1
timestamp 1700618825
transform 1 0 458 0 1 2168
box 231 427 920 2712
use 4T4R  x2
timestamp 1700618825
transform 1 0 458 0 1 -127
box 231 427 920 2712
use 4T4R  x3
timestamp 1700618825
transform 1 0 1154 0 1 2168
box 231 427 920 2712
use 4T4R  x4
timestamp 1700618825
transform 1 0 1154 0 1 -127
box 231 427 920 2712
<< labels >>
flabel metal2 689 3935 789 4035 0 FreeSans 128 0 0 0 WL1
port 0 nsew
flabel metal2 689 2779 789 2879 0 FreeSans 128 0 0 0 WL2
port 1 nsew
flabel metal2 689 1640 789 1740 0 FreeSans 128 0 0 0 WL3
port 2 nsew
flabel metal2 689 484 789 584 0 FreeSans 128 0 0 0 WL4
port 3 nsew
flabel metal3 1821 4780 1921 4880 0 FreeSans 128 0 0 0 SL4
port 11 nsew
flabel metal1 759 310 859 410 0 FreeSans 128 0 0 0 VSS
port 12 nsew
flabel metal3 778 4780 878 4880 0 FreeSans 128 0 0 0 SL1
port 8 nsew
flabel metal3 1474 4780 1574 4880 0 FreeSans 128 0 0 0 SL3
port 10 nsew
flabel metal3 1125 4780 1225 4880 0 FreeSans 128 0 0 0 SL2
port 9 nsew
flabel metal3 911 4780 1011 4880 0 FreeSans 128 0 0 0 BL1
port 4 nsew
flabel metal3 1258 4780 1358 4880 0 FreeSans 128 0 0 0 BL2
port 5 nsew
flabel metal3 1607 4780 1707 4880 0 FreeSans 128 0 0 0 BL3
port 6 nsew
flabel metal3 1954 4780 2054 4880 0 FreeSans 128 0 0 0 BL4
port 7 nsew
<< end >>
