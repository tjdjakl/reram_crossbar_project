magic
tech sky130B
magscale 1 2
timestamp 1700618825
<< metal1 >>
rect 4306 42240 4506 42440
rect 15578 40048 15778 40248
rect 12668 38820 12868 38846
rect 3250 38555 3450 38755
rect 12668 38660 12680 38820
rect 12860 38660 12870 38820
rect 12668 38646 12868 38660
rect 10414 38272 10614 38472
rect 2900 38000 3100 38200
rect 15578 31048 15778 31248
rect 12670 29660 12680 29820
rect 12860 29660 12870 29820
rect 2900 29000 3100 29200
rect 15578 22048 15778 22248
rect 12670 20660 12680 20820
rect 12860 20660 12870 20820
rect 2900 20000 3100 20200
rect 15578 13048 15778 13248
rect 12670 11660 12680 11820
rect 12860 11660 12870 11820
rect 2900 11000 3100 11200
rect 15578 4048 15778 4248
rect 12670 2660 12680 2820
rect 12860 2660 12870 2820
rect 2900 2000 3100 2200
rect 15578 -4952 15778 -4752
rect 12670 -6340 12680 -6180
rect 12860 -6340 12870 -6180
rect 2900 -7000 3100 -6800
rect 15578 -13952 15778 -13752
rect 12670 -15340 12680 -15180
rect 12860 -15340 12870 -15180
rect 2900 -16000 3100 -15800
rect 15579 -22952 15779 -22752
rect 12670 -24340 12680 -24180
rect 12860 -24340 12870 -24180
rect 2900 -25000 3100 -24800
<< via1 >>
rect 12680 38660 12860 38820
rect 12680 29660 12860 29820
rect 12680 20660 12860 20820
rect 12680 11660 12860 11820
rect 12680 2660 12860 2820
rect 12680 -6340 12860 -6180
rect 12680 -15340 12860 -15180
rect 12680 -24340 12860 -24180
<< metal2 >>
rect 13740 42520 13920 42530
rect 13740 42350 13920 42360
rect 12680 38820 12860 38830
rect 12680 38650 12860 38660
rect 13740 33500 13920 33510
rect 13740 33350 13920 33360
rect 12680 29820 12860 29830
rect 12680 29650 12860 29660
rect 13740 24500 13920 24510
rect 13740 24350 13920 24360
rect 12680 20820 12860 20830
rect 12680 20650 12860 20660
rect 13740 15500 13920 15510
rect 13740 15350 13920 15360
rect 12680 11820 12860 11830
rect 12680 11650 12860 11660
rect 13740 6500 13920 6510
rect 13740 6350 13920 6360
rect 12680 2820 12860 2830
rect 12680 2650 12860 2660
rect 13740 -2500 13920 -2490
rect 13740 -2650 13920 -2640
rect 12680 -6180 12860 -6170
rect 12680 -6350 12860 -6340
rect 13740 -11500 13920 -11490
rect 13740 -11650 13920 -11640
rect 12680 -15180 12860 -15170
rect 12680 -15350 12860 -15340
rect 13740 -20500 13920 -20490
rect 13740 -20650 13920 -20640
rect 12680 -24180 12860 -24170
rect 12680 -24350 12860 -24340
<< via2 >>
rect 13740 42360 13920 42520
rect 12680 38660 12860 38820
rect 13740 33360 13920 33500
rect 12680 29660 12860 29820
rect 13740 24360 13920 24500
rect 12680 20660 12860 20820
rect 13740 15360 13920 15500
rect 12680 11660 12860 11820
rect 13740 6360 13920 6500
rect 12680 2660 12860 2820
rect 13740 -2640 13920 -2500
rect 12680 -6340 12860 -6180
rect 13740 -11640 13920 -11500
rect 12680 -15340 12860 -15180
rect 13740 -20640 13920 -20500
rect 12680 -24340 12860 -24180
<< metal3 >>
rect 13730 42520 13930 42525
rect 13730 42360 13740 42520
rect 13920 42360 13930 42520
rect 13730 42355 13930 42360
rect 12670 38820 12870 38825
rect 3270 38580 3280 38720
rect 3420 38580 3430 38720
rect 12670 38660 12680 38820
rect 12860 38660 12870 38820
rect 12670 38655 12870 38660
rect 3250 29560 3260 29720
rect 3410 29560 3420 29720
rect 3270 20560 3280 20720
rect 3430 20560 3440 20720
rect 3270 11580 3280 11740
rect 3430 11580 3440 11740
rect 3270 2580 3280 2740
rect 3430 2580 3440 2740
rect 3270 -6420 3280 -6260
rect 3430 -6420 3440 -6260
rect 3270 -15420 3280 -15260
rect 3430 -15420 3440 -15260
rect 3270 -24420 3280 -24260
rect 3430 -24420 3440 -24260
rect 10440 -24660 10600 38380
rect 13740 33505 13920 42355
rect 13730 33500 13930 33505
rect 13730 33360 13740 33500
rect 13920 33360 13930 33500
rect 13730 33355 13930 33360
rect 12670 29820 12870 29825
rect 12670 29660 12680 29820
rect 12860 29660 12870 29820
rect 12670 29655 12870 29660
rect 12680 20825 12860 29655
rect 13740 24505 13920 33355
rect 13730 24500 13930 24505
rect 13730 24360 13740 24500
rect 13920 24360 13930 24500
rect 13730 24355 13930 24360
rect 12670 20820 12870 20825
rect 12670 20660 12680 20820
rect 12860 20660 12870 20820
rect 12670 20655 12870 20660
rect 12680 11825 12860 20655
rect 13740 15505 13920 24355
rect 13730 15500 13930 15505
rect 13730 15360 13740 15500
rect 13920 15360 13930 15500
rect 13730 15355 13930 15360
rect 12670 11820 12870 11825
rect 12670 11660 12680 11820
rect 12860 11660 12870 11820
rect 12670 11655 12870 11660
rect 12680 2825 12860 11655
rect 13740 6505 13920 15355
rect 13730 6500 13930 6505
rect 13730 6360 13740 6500
rect 13920 6360 13930 6500
rect 13730 6355 13930 6360
rect 12670 2820 12870 2825
rect 12670 2660 12680 2820
rect 12860 2660 12870 2820
rect 12670 2655 12870 2660
rect 12680 -6175 12860 2655
rect 13740 -2495 13920 6355
rect 13730 -2500 13930 -2495
rect 13730 -2640 13740 -2500
rect 13920 -2640 13930 -2500
rect 13730 -2645 13930 -2640
rect 12670 -6180 12870 -6175
rect 12670 -6340 12680 -6180
rect 12860 -6340 12870 -6180
rect 12670 -6345 12870 -6340
rect 12680 -15175 12860 -6345
rect 13740 -11495 13920 -2645
rect 13730 -11500 13930 -11495
rect 13730 -11640 13740 -11500
rect 13920 -11640 13930 -11500
rect 13730 -11645 13930 -11640
rect 12670 -15180 12870 -15175
rect 12670 -15340 12680 -15180
rect 12860 -15340 12870 -15180
rect 12670 -15345 12870 -15340
rect 12680 -24175 12860 -15345
rect 13740 -20495 13920 -11645
rect 13730 -20500 13930 -20495
rect 13730 -20640 13740 -20500
rect 13920 -20640 13930 -20500
rect 13730 -20645 13930 -20640
rect 12670 -24180 12870 -24175
rect 12670 -24340 12680 -24180
rect 12860 -24340 12870 -24180
rect 12670 -24345 12870 -24340
<< via3 >>
rect 3280 38580 3420 38720
rect 3260 29560 3410 29720
rect 3280 20560 3430 20720
rect 3280 11580 3430 11740
rect 3280 2580 3430 2740
rect 3280 -6420 3430 -6260
rect 3280 -15420 3430 -15260
rect 3280 -24420 3430 -24260
<< metal4 >>
rect 3279 38720 3421 38721
rect 3279 38580 3280 38720
rect 3420 38580 3421 38720
rect 3279 38579 3421 38580
rect 3280 29721 3420 38579
rect 3259 29720 3420 29721
rect 3259 29560 3260 29720
rect 3410 29560 3420 29720
rect 3259 29559 3420 29560
rect 3280 20721 3420 29559
rect 3279 20720 3431 20721
rect 3279 20560 3280 20720
rect 3430 20560 3431 20720
rect 3279 20559 3431 20560
rect 3280 11741 3420 20559
rect 3279 11740 3431 11741
rect 3279 11580 3280 11740
rect 3430 11580 3431 11740
rect 3279 11579 3431 11580
rect 3280 2741 3420 11579
rect 3279 2740 3431 2741
rect 3279 2580 3280 2740
rect 3430 2580 3431 2740
rect 3279 2579 3431 2580
rect 3280 -6259 3420 2579
rect 3279 -6260 3431 -6259
rect 3279 -6420 3280 -6260
rect 3430 -6420 3431 -6260
rect 3279 -6421 3431 -6420
rect 3280 -15259 3420 -6421
rect 3279 -15260 3431 -15259
rect 3279 -15420 3280 -15260
rect 3430 -15420 3431 -15260
rect 3279 -15421 3431 -15420
rect 3280 -24259 3420 -15421
rect 3279 -24260 3431 -24259
rect 3279 -24420 3280 -24260
rect 3430 -24420 3431 -24260
rect 3279 -24421 3431 -24420
use 1LineSelectOutput04  x1
timestamp 1700618825
transform 1 0 -752 0 1 37496
box 3752 504 16530 9374
use 1LineSelectOutput04  x2
timestamp 1700618825
transform 1 0 -752 0 1 28496
box 3752 504 16530 9374
use 1LineSelectOutput04  x3
timestamp 1700618825
transform 1 0 -752 0 1 19496
box 3752 504 16530 9374
use 1LineSelectOutput04  x4
timestamp 1700618825
transform 1 0 -752 0 1 10496
box 3752 504 16530 9374
use 1LineSelectOutput04  x5
timestamp 1700618825
transform 1 0 -752 0 1 1496
box 3752 504 16530 9374
use 1LineSelectOutput04  x6
timestamp 1700618825
transform 1 0 -752 0 1 -7504
box 3752 504 16530 9374
use 1LineSelectOutput04  x7
timestamp 1700618825
transform 1 0 -752 0 1 -16504
box 3752 504 16530 9374
use 1LineSelectOutput04  x8
timestamp 1700618825
transform 1 0 -752 0 1 -25504
box 3752 504 16530 9374
<< labels >>
flabel metal1 10414 38272 10614 38472 0 FreeSans 256 0 0 0 Gnd
port 20 nsew
flabel metal1 15579 -22952 15779 -22752 0 FreeSans 256 0 0 0 LA_OUT8
port 19 nsew
flabel metal1 15578 -13952 15778 -13752 0 FreeSans 256 0 0 0 LA_OUT7
port 18 nsew
flabel metal1 15578 -4952 15778 -4752 0 FreeSans 256 0 0 0 LA_OUT6
port 17 nsew
flabel metal1 15578 4048 15778 4248 0 FreeSans 256 0 0 0 LA_OUT5
port 16 nsew
flabel metal1 15578 13048 15778 13248 0 FreeSans 256 0 0 0 LA_OUT4
port 15 nsew
flabel metal1 15578 22048 15778 22248 0 FreeSans 256 0 0 0 LA_OUT3
port 14 nsew
flabel metal1 15578 31048 15778 31248 0 FreeSans 256 0 0 0 LA_OUT2
port 13 nsew
flabel metal1 15578 40048 15778 40248 0 FreeSans 256 0 0 0 LA_OUT1
port 12 nsew
flabel metal1 3250 38555 3450 38755 0 FreeSans 256 0 0 0 VSSneg
port 11 nsew
flabel metal1 12668 38646 12868 38846 0 FreeSans 256 0 0 0 VSS
port 10 nsew
flabel metal1 4306 42240 4506 42440 0 FreeSans 256 0 0 0 VDD18
port 9 nsew
flabel metal1 2900 38000 3100 38200 0 FreeSans 256 0 0 0 SL_LA_OUT1
port 0 nsew
flabel metal1 2900 -25000 3100 -24800 0 FreeSans 256 0 0 0 SL_LA_OUT8
port 8 nsew
flabel metal1 2900 -16000 3100 -15800 0 FreeSans 256 0 0 0 SL_LA_OUT7
port 7 nsew
flabel metal1 2900 -7000 3100 -6800 0 FreeSans 256 0 0 0 SL_LA_OUT6
port 5 nsew
flabel metal1 2900 2000 3100 2200 0 FreeSans 256 0 0 0 SL_LA_OUT5
port 4 nsew
flabel metal1 2900 11000 3100 11200 0 FreeSans 256 0 0 0 SL_LA_OUT4
port 3 nsew
flabel metal1 2900 20000 3100 20200 0 FreeSans 256 0 0 0 SL_LA_OUT3
port 2 nsew
flabel metal1 2900 29000 3100 29200 0 FreeSans 256 0 0 0 SL_LA_OUT2
port 1 nsew
<< end >>
