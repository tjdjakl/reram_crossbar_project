magic
tech sky130B
magscale 1 2
timestamp 1700618825
<< metal1 >>
rect 91617 88543 91817 88743
rect 102890 86352 103090 86552
rect 99980 85120 100180 85149
rect 90554 84860 90754 85060
rect 99980 84960 100000 85120
rect 100160 84960 100180 85120
rect 99980 84949 100180 84960
rect 90300 84400 90500 84600
rect 97725 84576 97925 84776
rect 102889 74352 103089 74552
rect 99990 72980 100000 73140
rect 100160 72980 100170 73140
rect 90300 72400 90500 72600
rect 102890 62353 103090 62553
rect 99990 60980 100000 61140
rect 100160 60980 100170 61140
rect 90300 60400 90500 60600
rect 102890 50352 103090 50552
rect 99990 48980 100000 49140
rect 100160 48980 100170 49140
rect 90300 48400 90500 48600
rect 102889 38352 103089 38552
rect 99990 36980 100000 37140
rect 100160 36980 100170 37140
rect 90300 36400 90500 36600
rect 102890 26352 103090 26552
rect 99990 24980 100000 25140
rect 100160 24980 100170 25140
rect 90300 24400 90500 24600
rect 102890 14352 103090 14552
rect 99990 12980 100000 13140
rect 100160 12980 100170 13140
rect 90300 12400 90500 12600
rect 102890 2352 103090 2552
rect 99990 980 100000 1140
rect 100160 980 100170 1140
rect 90300 400 90500 600
<< via1 >>
rect 100000 84960 100160 85120
rect 100000 72980 100160 73140
rect 100000 60980 100160 61140
rect 100000 48980 100160 49140
rect 100000 36980 100160 37140
rect 100000 24980 100160 25140
rect 100000 12980 100160 13140
rect 100000 980 100160 1140
<< metal2 >>
rect 101060 88800 101220 88810
rect 101060 88650 101220 88660
rect 100000 85120 100160 85130
rect 100000 84950 100160 84960
rect 101060 76800 101220 76810
rect 101060 76650 101220 76660
rect 100000 73140 100160 73150
rect 100000 72970 100160 72980
rect 101060 64800 101220 64810
rect 101060 64650 101220 64660
rect 100000 61140 100160 61150
rect 100000 60970 100160 60980
rect 101060 52800 101220 52810
rect 101060 52650 101220 52660
rect 100000 49140 100160 49150
rect 100000 48970 100160 48980
rect 101060 40800 101220 40810
rect 101060 40650 101220 40660
rect 100000 37140 100160 37150
rect 100000 36970 100160 36980
rect 101060 28800 101220 28810
rect 101060 28650 101220 28660
rect 100000 25140 100160 25150
rect 100000 24970 100160 24980
rect 101060 16800 101220 16810
rect 101060 16650 101220 16660
rect 100000 13140 100160 13150
rect 100000 12970 100160 12980
rect 101060 4800 101220 4810
rect 101060 4650 101220 4660
rect 100000 1140 100160 1150
rect 100000 970 100160 980
<< via2 >>
rect 101060 88660 101220 88800
rect 100000 84960 100160 85120
rect 101060 76660 101220 76800
rect 100000 72980 100160 73140
rect 101060 64660 101220 64800
rect 100000 60980 100160 61140
rect 101060 52660 101220 52800
rect 100000 48980 100160 49140
rect 101060 40660 101220 40800
rect 100000 36980 100160 37140
rect 101060 28660 101220 28800
rect 100000 24980 100160 25140
rect 101060 16660 101220 16800
rect 100000 12980 100160 13140
rect 101060 4660 101220 4800
rect 100000 980 100160 1140
<< metal3 >>
rect 101050 88800 101230 88805
rect 101050 88660 101060 88800
rect 101220 88660 101230 88800
rect 101050 88655 101230 88660
rect 99990 85120 100170 85125
rect 90570 84880 90580 85040
rect 90740 84880 90750 85040
rect 99990 84960 100000 85120
rect 100160 84960 100170 85120
rect 99990 84955 100170 84960
rect 90570 72880 90580 73040
rect 90740 72880 90750 73040
rect 90570 60880 90580 61040
rect 90740 60880 90750 61040
rect 90570 48880 90580 49040
rect 90740 48880 90750 49040
rect 90570 36880 90580 37040
rect 90740 36880 90750 37040
rect 90570 24880 90580 25040
rect 90740 24880 90750 25040
rect 90570 12880 90580 13040
rect 90740 12880 90750 13040
rect 90570 880 90580 1040
rect 90740 880 90750 1040
rect 97740 660 97900 84660
rect 100000 73145 100160 84955
rect 101060 76805 101220 88655
rect 101050 76800 101230 76805
rect 101050 76660 101060 76800
rect 101220 76660 101230 76800
rect 101050 76655 101230 76660
rect 99990 73140 100170 73145
rect 99990 72980 100000 73140
rect 100160 72980 100170 73140
rect 99990 72975 100170 72980
rect 100000 61145 100160 72975
rect 101060 64805 101220 76655
rect 101050 64800 101230 64805
rect 101050 64660 101060 64800
rect 101220 64660 101230 64800
rect 101050 64655 101230 64660
rect 99990 61140 100170 61145
rect 99990 60980 100000 61140
rect 100160 60980 100170 61140
rect 99990 60975 100170 60980
rect 100000 49145 100160 60975
rect 101060 52805 101220 64655
rect 101050 52800 101230 52805
rect 101050 52660 101060 52800
rect 101220 52660 101230 52800
rect 101050 52655 101230 52660
rect 99990 49140 100170 49145
rect 99990 48980 100000 49140
rect 100160 48980 100170 49140
rect 99990 48975 100170 48980
rect 100000 37145 100160 48975
rect 101060 40805 101220 52655
rect 101050 40800 101230 40805
rect 101050 40660 101060 40800
rect 101220 40660 101230 40800
rect 101050 40655 101230 40660
rect 99990 37140 100170 37145
rect 99990 36980 100000 37140
rect 100160 36980 100170 37140
rect 99990 36975 100170 36980
rect 100000 25145 100160 36975
rect 101060 28805 101220 40655
rect 101050 28800 101230 28805
rect 101050 28660 101060 28800
rect 101220 28660 101230 28800
rect 101050 28655 101230 28660
rect 99990 25140 100170 25145
rect 99990 24980 100000 25140
rect 100160 24980 100170 25140
rect 99990 24975 100170 24980
rect 100000 13145 100160 24975
rect 101060 16805 101220 28655
rect 101050 16800 101230 16805
rect 101050 16660 101060 16800
rect 101220 16660 101230 16800
rect 101050 16655 101230 16660
rect 99990 13140 100170 13145
rect 99990 12980 100000 13140
rect 100160 12980 100170 13140
rect 99990 12975 100170 12980
rect 100000 1145 100160 12975
rect 101060 4805 101220 16655
rect 101050 4800 101230 4805
rect 101050 4660 101060 4800
rect 101220 4660 101230 4800
rect 101050 4655 101230 4660
rect 99990 1140 100170 1145
rect 99990 980 100000 1140
rect 100160 980 100170 1140
rect 99990 975 100170 980
<< via3 >>
rect 90580 84880 90740 85040
rect 90580 72880 90740 73040
rect 90580 60880 90740 61040
rect 90580 48880 90740 49040
rect 90580 36880 90740 37040
rect 90580 24880 90740 25040
rect 90580 12880 90740 13040
rect 90580 880 90740 1040
<< metal4 >>
rect 90579 85040 90741 85041
rect 90579 84880 90580 85040
rect 90740 84880 90741 85040
rect 90579 84879 90741 84880
rect 90580 73041 90740 84879
rect 90579 73040 90741 73041
rect 90579 72880 90580 73040
rect 90740 72880 90741 73040
rect 90579 72879 90741 72880
rect 90580 61041 90740 72879
rect 90579 61040 90741 61041
rect 90579 60880 90580 61040
rect 90740 60880 90741 61040
rect 90579 60879 90741 60880
rect 90580 49041 90740 60879
rect 90579 49040 90741 49041
rect 90579 48880 90580 49040
rect 90740 48880 90741 49040
rect 90579 48879 90741 48880
rect 90580 37041 90740 48879
rect 90579 37040 90741 37041
rect 90579 36880 90580 37040
rect 90740 36880 90741 37040
rect 90579 36879 90741 36880
rect 90580 25041 90740 36879
rect 90579 25040 90741 25041
rect 90579 24880 90580 25040
rect 90740 24880 90741 25040
rect 90579 24879 90741 24880
rect 90580 13041 90740 24879
rect 90579 13040 90741 13041
rect 90579 12880 90580 13040
rect 90740 12880 90741 13040
rect 90579 12879 90741 12880
rect 90580 1041 90740 12879
rect 90579 1040 90741 1041
rect 90579 880 90580 1040
rect 90740 880 90741 1040
rect 90579 879 90741 880
use 1LineSelectOutput02  x1
timestamp 1700618825
transform 1 0 86560 0 1 83800
box 3640 600 16530 12482
use 1LineSelectOutput02  x2
timestamp 1700618825
transform 1 0 86560 0 1 71800
box 3640 600 16530 12482
use 1LineSelectOutput02  x3
timestamp 1700618825
transform 1 0 86560 0 1 59800
box 3640 600 16530 12482
use 1LineSelectOutput02  x4
timestamp 1700618825
transform 1 0 86560 0 1 47800
box 3640 600 16530 12482
use 1LineSelectOutput02  x5
timestamp 1700618825
transform 1 0 86560 0 1 35800
box 3640 600 16530 12482
use 1LineSelectOutput02  x6
timestamp 1700618825
transform 1 0 86560 0 1 23800
box 3640 600 16530 12482
use 1LineSelectOutput02  x7
timestamp 1700618825
transform 1 0 86560 0 1 11800
box 3640 600 16530 12482
use 1LineSelectOutput02  x8
timestamp 1700618825
transform 1 0 86560 0 1 -200
box 3640 600 16530 12482
<< labels >>
flabel metal1 90300 84400 90500 84600 0 FreeSans 256 0 0 0 SL_LA_OUT1
port 0 nsew
flabel metal1 90300 72400 90500 72600 0 FreeSans 256 0 0 0 SL_LA_OUT2
port 1 nsew
flabel metal1 90300 60400 90500 60600 0 FreeSans 256 0 0 0 SL_LA_OUT3
port 2 nsew
flabel metal1 90300 48400 90500 48600 0 FreeSans 256 0 0 0 SL_LA_OUT4
port 3 nsew
flabel metal1 90300 36400 90500 36600 0 FreeSans 256 0 0 0 SL_LA_OUT5
port 4 nsew
flabel metal1 90300 24400 90500 24600 0 FreeSans 256 0 0 0 SL_LA_OUT6
port 5 nsew
flabel metal1 90300 12400 90500 12600 0 FreeSans 256 0 0 0 SL_LA_OUT7
port 7 nsew
flabel metal1 90300 400 90500 600 0 FreeSans 256 0 0 0 SL_LA_OUT8
port 8 nsew
flabel metal1 91617 88543 91817 88743 0 FreeSans 256 0 0 0 VDD18
port 9 nsew
flabel metal1 99980 84949 100180 85149 0 FreeSans 256 0 0 0 VSS
port 10 nsew
flabel metal1 90554 84860 90754 85060 0 FreeSans 256 0 0 0 VSSneg
port 11 nsew
flabel metal1 97725 84576 97925 84776 0 FreeSans 256 0 0 0 Gnd
port 20 nsew
flabel metal1 102890 86352 103090 86552 0 FreeSans 256 0 0 0 LA_OUT1
port 12 nsew
flabel metal1 102889 74352 103089 74552 0 FreeSans 256 0 0 0 LA_OUT2
port 13 nsew
flabel metal1 102890 62353 103090 62553 0 FreeSans 256 0 0 0 LA_OUT3
port 14 nsew
flabel metal1 102890 50352 103090 50552 0 FreeSans 256 0 0 0 LA_OUT4
port 15 nsew
flabel metal1 102889 38352 103089 38552 0 FreeSans 256 0 0 0 LA_OUT5
port 16 nsew
flabel metal1 102890 26352 103090 26552 0 FreeSans 256 0 0 0 LA_OUT6
port 17 nsew
flabel metal1 102890 14352 103090 14552 0 FreeSans 256 0 0 0 LA_OUT7
port 18 nsew
flabel metal1 102890 2352 103090 2552 0 FreeSans 256 0 0 0 LA_OUT8
port 19 nsew
<< end >>
