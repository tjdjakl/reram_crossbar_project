magic
tech sky130B
magscale 1 2
timestamp 1688980957
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808615  sky130_fd_pr__model__nfet_highvoltage__example_55959141808615_0
timestamp 1688980957
transform 1 0 119 0 -1 284
box -1 0 649 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808616  sky130_fd_pr__model__pfet_highvoltage__example_55959141808616_0
timestamp 1688980957
transform 1 0 119 0 -1 682
box -1 0 649 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808616  sky130_fd_pr__model__pfet_highvoltage__example_55959141808616_1
timestamp 1688980957
transform 1 0 119 0 1 750
box -1 0 649 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1688980957
transform 0 -1 812 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1688980957
transform 0 -1 812 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1688980957
transform 0 -1 108 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1688980957
transform 0 -1 460 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1688980957
transform 0 -1 460 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1688980957
transform 0 -1 108 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1688980957
transform 0 -1 215 1 0 316
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1688980957
transform 0 -1 737 1 0 316
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808612  sky130_fd_pr__via_pol1__example_55959141808612_0
timestamp 1688980957
transform 1 0 302 0 1 341
box 0 0 1 1
<< properties >>
string GDS_END 7954714
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7950372
<< end >>
