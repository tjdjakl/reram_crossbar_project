magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< dnwell >>
rect 640 9736 14336 36182
<< nwell >>
rect 531 35918 14447 36293
rect 531 10000 846 35918
rect 14072 10000 14447 35918
rect 531 9569 14447 10000
<< pwell >>
rect 219 36363 14750 36600
rect 219 9554 456 36363
rect 1151 34538 13843 34710
rect 1151 10360 1323 34538
rect 13671 10360 13843 34538
rect 1151 10188 13843 10360
rect 14513 9554 14750 36363
rect 219 9317 14750 9554
<< mvpsubdiff >>
rect 245 36499 14724 36574
rect 245 36465 492 36499
rect 526 36465 560 36499
rect 594 36465 628 36499
rect 662 36465 696 36499
rect 730 36465 764 36499
rect 798 36465 832 36499
rect 866 36465 900 36499
rect 934 36465 968 36499
rect 1002 36465 1036 36499
rect 1070 36465 1104 36499
rect 1138 36465 1172 36499
rect 1206 36465 1240 36499
rect 1274 36465 1308 36499
rect 1342 36465 1376 36499
rect 1410 36465 1444 36499
rect 1478 36465 1512 36499
rect 1546 36465 1580 36499
rect 1614 36465 1648 36499
rect 1682 36465 1716 36499
rect 1750 36465 1784 36499
rect 1818 36465 1852 36499
rect 1886 36465 1920 36499
rect 1954 36465 1988 36499
rect 2022 36465 2056 36499
rect 2090 36465 2124 36499
rect 2158 36465 2192 36499
rect 2226 36465 2260 36499
rect 2294 36465 2328 36499
rect 2362 36465 2396 36499
rect 2430 36465 2464 36499
rect 2498 36465 2532 36499
rect 2566 36465 2600 36499
rect 2634 36465 2668 36499
rect 2702 36465 2736 36499
rect 2770 36465 2804 36499
rect 2838 36465 2872 36499
rect 2906 36465 2940 36499
rect 2974 36465 3008 36499
rect 3042 36465 3076 36499
rect 3110 36465 3144 36499
rect 3178 36465 3212 36499
rect 3246 36465 3280 36499
rect 3314 36465 3348 36499
rect 3382 36465 3416 36499
rect 3450 36465 3484 36499
rect 3518 36465 3552 36499
rect 3586 36465 3620 36499
rect 3654 36465 3688 36499
rect 3722 36465 3756 36499
rect 3790 36465 3824 36499
rect 3858 36465 3892 36499
rect 3926 36465 3960 36499
rect 3994 36465 4028 36499
rect 4062 36465 4096 36499
rect 4130 36465 4164 36499
rect 4198 36465 4232 36499
rect 4266 36465 4300 36499
rect 4334 36465 4368 36499
rect 4402 36465 4436 36499
rect 4470 36465 4504 36499
rect 4538 36465 4572 36499
rect 4606 36465 4640 36499
rect 4674 36465 4708 36499
rect 4742 36465 4776 36499
rect 4810 36465 4844 36499
rect 4878 36465 4912 36499
rect 4946 36465 4980 36499
rect 5014 36465 5048 36499
rect 5082 36465 5116 36499
rect 5150 36465 5184 36499
rect 5218 36465 5252 36499
rect 5286 36465 5320 36499
rect 5354 36465 5388 36499
rect 5422 36465 5456 36499
rect 5490 36465 5524 36499
rect 5558 36465 5592 36499
rect 5626 36465 5660 36499
rect 5694 36465 5728 36499
rect 5762 36465 5796 36499
rect 5830 36465 5864 36499
rect 5898 36465 5932 36499
rect 5966 36465 6000 36499
rect 6034 36465 6068 36499
rect 6102 36465 6136 36499
rect 6170 36465 6204 36499
rect 6238 36465 6272 36499
rect 6306 36465 6340 36499
rect 6374 36465 6408 36499
rect 6442 36465 6476 36499
rect 6510 36465 6544 36499
rect 6578 36465 6612 36499
rect 6646 36465 6680 36499
rect 6714 36465 6748 36499
rect 6782 36465 6816 36499
rect 6850 36465 6884 36499
rect 6918 36465 6952 36499
rect 6986 36465 7020 36499
rect 7054 36465 7088 36499
rect 7122 36465 7156 36499
rect 7190 36465 7224 36499
rect 7258 36465 7292 36499
rect 7326 36465 7360 36499
rect 7394 36465 7428 36499
rect 7462 36465 7496 36499
rect 7530 36465 7564 36499
rect 7598 36465 7632 36499
rect 7666 36465 7700 36499
rect 7734 36465 7768 36499
rect 7802 36465 7836 36499
rect 7870 36465 7904 36499
rect 7938 36465 7972 36499
rect 8006 36465 8040 36499
rect 8074 36465 8108 36499
rect 8142 36465 8176 36499
rect 8210 36465 8244 36499
rect 8278 36465 8312 36499
rect 8346 36465 8380 36499
rect 8414 36465 8448 36499
rect 8482 36465 8516 36499
rect 8550 36465 8584 36499
rect 8618 36465 8652 36499
rect 8686 36465 8720 36499
rect 8754 36465 8788 36499
rect 8822 36465 8856 36499
rect 8890 36465 8924 36499
rect 8958 36465 8992 36499
rect 9026 36465 9060 36499
rect 9094 36465 9128 36499
rect 9162 36465 9196 36499
rect 9230 36465 9264 36499
rect 9298 36465 9332 36499
rect 9366 36465 9400 36499
rect 9434 36465 9468 36499
rect 9502 36465 9536 36499
rect 9570 36465 9604 36499
rect 9638 36465 9672 36499
rect 9706 36465 9740 36499
rect 9774 36465 9808 36499
rect 9842 36465 9876 36499
rect 9910 36465 9944 36499
rect 9978 36465 10012 36499
rect 10046 36465 10080 36499
rect 10114 36465 10148 36499
rect 10182 36465 10216 36499
rect 10250 36465 10284 36499
rect 10318 36465 10352 36499
rect 10386 36465 10420 36499
rect 10454 36465 10488 36499
rect 10522 36465 10556 36499
rect 10590 36465 10624 36499
rect 10658 36465 10692 36499
rect 10726 36465 10760 36499
rect 10794 36465 10828 36499
rect 10862 36465 10896 36499
rect 10930 36465 10964 36499
rect 10998 36465 11032 36499
rect 11066 36465 11100 36499
rect 11134 36465 11168 36499
rect 11202 36465 11236 36499
rect 11270 36465 11304 36499
rect 11338 36465 11372 36499
rect 11406 36465 11440 36499
rect 11474 36465 11508 36499
rect 11542 36465 11576 36499
rect 11610 36465 11644 36499
rect 11678 36465 11712 36499
rect 11746 36465 11780 36499
rect 11814 36465 11848 36499
rect 11882 36465 11916 36499
rect 11950 36465 11984 36499
rect 12018 36465 12052 36499
rect 12086 36465 12120 36499
rect 12154 36465 12188 36499
rect 12222 36465 12256 36499
rect 12290 36465 12324 36499
rect 12358 36465 12392 36499
rect 12426 36465 12460 36499
rect 12494 36465 12528 36499
rect 12562 36465 12596 36499
rect 12630 36465 12664 36499
rect 12698 36465 12732 36499
rect 12766 36465 12800 36499
rect 12834 36465 12868 36499
rect 12902 36465 12936 36499
rect 12970 36465 13004 36499
rect 13038 36465 13072 36499
rect 13106 36465 13140 36499
rect 13174 36465 13208 36499
rect 13242 36465 13276 36499
rect 13310 36465 13344 36499
rect 13378 36465 13412 36499
rect 13446 36465 13480 36499
rect 13514 36465 13548 36499
rect 13582 36465 13616 36499
rect 13650 36465 13684 36499
rect 13718 36465 13752 36499
rect 13786 36465 13820 36499
rect 13854 36465 13888 36499
rect 13922 36465 13956 36499
rect 13990 36465 14024 36499
rect 14058 36465 14092 36499
rect 14126 36465 14160 36499
rect 14194 36465 14228 36499
rect 14262 36465 14296 36499
rect 14330 36465 14364 36499
rect 14398 36465 14432 36499
rect 14466 36465 14724 36499
rect 245 36389 14724 36465
rect 245 36335 430 36389
rect 245 36301 322 36335
rect 356 36301 430 36335
rect 245 36267 430 36301
rect 245 36233 322 36267
rect 356 36233 430 36267
rect 245 36199 430 36233
rect 14539 36327 14724 36389
rect 14539 36293 14609 36327
rect 14643 36293 14724 36327
rect 14539 36259 14724 36293
rect 245 36165 322 36199
rect 356 36165 430 36199
rect 245 36131 430 36165
rect 245 36097 322 36131
rect 356 36097 430 36131
rect 245 36063 430 36097
rect 245 36029 322 36063
rect 356 36029 430 36063
rect 245 35995 430 36029
rect 245 35961 322 35995
rect 356 35961 430 35995
rect 245 35927 430 35961
rect 245 35893 322 35927
rect 356 35893 430 35927
rect 245 35859 430 35893
rect 245 35825 322 35859
rect 356 35825 430 35859
rect 245 35791 430 35825
rect 245 35757 322 35791
rect 356 35757 430 35791
rect 245 35723 430 35757
rect 245 35689 322 35723
rect 356 35689 430 35723
rect 245 35655 430 35689
rect 245 35621 322 35655
rect 356 35621 430 35655
rect 245 35587 430 35621
rect 245 35553 322 35587
rect 356 35553 430 35587
rect 245 35519 430 35553
rect 245 35485 322 35519
rect 356 35485 430 35519
rect 245 35451 430 35485
rect 245 35417 322 35451
rect 356 35417 430 35451
rect 245 35383 430 35417
rect 245 35349 322 35383
rect 356 35349 430 35383
rect 245 35315 430 35349
rect 245 35281 322 35315
rect 356 35281 430 35315
rect 245 35247 430 35281
rect 245 35213 322 35247
rect 356 35213 430 35247
rect 245 35179 430 35213
rect 245 35145 322 35179
rect 356 35145 430 35179
rect 245 35111 430 35145
rect 245 35077 322 35111
rect 356 35077 430 35111
rect 245 35043 430 35077
rect 245 35009 322 35043
rect 356 35009 430 35043
rect 245 34975 430 35009
rect 245 34941 322 34975
rect 356 34941 430 34975
rect 245 34907 430 34941
rect 245 34873 322 34907
rect 356 34873 430 34907
rect 245 34839 430 34873
rect 245 34805 322 34839
rect 356 34805 430 34839
rect 245 34771 430 34805
rect 245 34737 322 34771
rect 356 34737 430 34771
rect 245 34703 430 34737
rect 245 34669 322 34703
rect 356 34669 430 34703
rect 245 34635 430 34669
rect 245 34601 322 34635
rect 356 34601 430 34635
rect 245 34567 430 34601
rect 245 34533 322 34567
rect 356 34533 430 34567
rect 245 34499 430 34533
rect 245 34465 322 34499
rect 356 34465 430 34499
rect 245 34431 430 34465
rect 245 34397 322 34431
rect 356 34397 430 34431
rect 245 34363 430 34397
rect 245 34329 322 34363
rect 356 34329 430 34363
rect 245 34295 430 34329
rect 245 34261 322 34295
rect 356 34261 430 34295
rect 245 34227 430 34261
rect 245 34193 322 34227
rect 356 34193 430 34227
rect 245 34159 430 34193
rect 245 34125 322 34159
rect 356 34125 430 34159
rect 245 34091 430 34125
rect 245 34057 322 34091
rect 356 34057 430 34091
rect 245 34023 430 34057
rect 245 33989 322 34023
rect 356 33989 430 34023
rect 245 33955 430 33989
rect 245 33921 322 33955
rect 356 33921 430 33955
rect 245 33887 430 33921
rect 245 33853 322 33887
rect 356 33853 430 33887
rect 245 33819 430 33853
rect 245 33785 322 33819
rect 356 33785 430 33819
rect 245 33751 430 33785
rect 245 33717 322 33751
rect 356 33717 430 33751
rect 245 33683 430 33717
rect 245 33649 322 33683
rect 356 33649 430 33683
rect 245 33615 430 33649
rect 245 33581 322 33615
rect 356 33581 430 33615
rect 245 33547 430 33581
rect 245 33513 322 33547
rect 356 33513 430 33547
rect 245 33479 430 33513
rect 245 33445 322 33479
rect 356 33445 430 33479
rect 245 33411 430 33445
rect 245 33377 322 33411
rect 356 33377 430 33411
rect 245 33343 430 33377
rect 245 33309 322 33343
rect 356 33309 430 33343
rect 245 33275 430 33309
rect 245 33241 322 33275
rect 356 33241 430 33275
rect 245 33207 430 33241
rect 245 33173 322 33207
rect 356 33173 430 33207
rect 245 33139 430 33173
rect 245 33105 322 33139
rect 356 33105 430 33139
rect 245 33071 430 33105
rect 245 33037 322 33071
rect 356 33037 430 33071
rect 245 33003 430 33037
rect 245 32969 322 33003
rect 356 32969 430 33003
rect 245 32935 430 32969
rect 245 32901 322 32935
rect 356 32901 430 32935
rect 245 32867 430 32901
rect 245 32833 322 32867
rect 356 32833 430 32867
rect 245 32799 430 32833
rect 245 32765 322 32799
rect 356 32765 430 32799
rect 245 32731 430 32765
rect 245 32697 322 32731
rect 356 32697 430 32731
rect 245 32663 430 32697
rect 245 32629 322 32663
rect 356 32629 430 32663
rect 245 32595 430 32629
rect 245 32561 322 32595
rect 356 32561 430 32595
rect 245 32527 430 32561
rect 245 32493 322 32527
rect 356 32493 430 32527
rect 245 32459 430 32493
rect 245 32425 322 32459
rect 356 32425 430 32459
rect 245 32391 430 32425
rect 245 32357 322 32391
rect 356 32357 430 32391
rect 245 32323 430 32357
rect 245 32289 322 32323
rect 356 32289 430 32323
rect 245 32255 430 32289
rect 245 32221 322 32255
rect 356 32221 430 32255
rect 245 32187 430 32221
rect 245 32153 322 32187
rect 356 32153 430 32187
rect 245 32119 430 32153
rect 245 32085 322 32119
rect 356 32085 430 32119
rect 245 32051 430 32085
rect 245 32017 322 32051
rect 356 32017 430 32051
rect 245 31983 430 32017
rect 245 31949 322 31983
rect 356 31949 430 31983
rect 245 31915 430 31949
rect 245 31881 322 31915
rect 356 31881 430 31915
rect 245 31847 430 31881
rect 245 31813 322 31847
rect 356 31813 430 31847
rect 245 31779 430 31813
rect 245 31745 322 31779
rect 356 31745 430 31779
rect 245 31711 430 31745
rect 245 31677 322 31711
rect 356 31677 430 31711
rect 245 31643 430 31677
rect 245 31609 322 31643
rect 356 31609 430 31643
rect 245 31575 430 31609
rect 245 31541 322 31575
rect 356 31541 430 31575
rect 245 31507 430 31541
rect 245 31473 322 31507
rect 356 31473 430 31507
rect 245 31439 430 31473
rect 245 31405 322 31439
rect 356 31405 430 31439
rect 245 31371 430 31405
rect 245 31337 322 31371
rect 356 31337 430 31371
rect 245 31303 430 31337
rect 245 31269 322 31303
rect 356 31269 430 31303
rect 245 31235 430 31269
rect 245 31201 322 31235
rect 356 31201 430 31235
rect 245 31167 430 31201
rect 245 31133 322 31167
rect 356 31133 430 31167
rect 245 31099 430 31133
rect 245 31065 322 31099
rect 356 31065 430 31099
rect 245 31031 430 31065
rect 245 30997 322 31031
rect 356 30997 430 31031
rect 245 30963 430 30997
rect 245 30929 322 30963
rect 356 30929 430 30963
rect 245 30895 430 30929
rect 245 30861 322 30895
rect 356 30861 430 30895
rect 245 30827 430 30861
rect 245 30793 322 30827
rect 356 30793 430 30827
rect 245 30759 430 30793
rect 245 30725 322 30759
rect 356 30725 430 30759
rect 245 30691 430 30725
rect 245 30657 322 30691
rect 356 30657 430 30691
rect 245 30623 430 30657
rect 245 30589 322 30623
rect 356 30589 430 30623
rect 245 30555 430 30589
rect 245 30521 322 30555
rect 356 30521 430 30555
rect 245 30487 430 30521
rect 245 30453 322 30487
rect 356 30453 430 30487
rect 245 30419 430 30453
rect 245 30385 322 30419
rect 356 30385 430 30419
rect 245 30351 430 30385
rect 245 30317 322 30351
rect 356 30317 430 30351
rect 245 30283 430 30317
rect 245 30249 322 30283
rect 356 30249 430 30283
rect 245 30215 430 30249
rect 245 30181 322 30215
rect 356 30181 430 30215
rect 245 30147 430 30181
rect 245 30113 322 30147
rect 356 30113 430 30147
rect 245 30079 430 30113
rect 245 30045 322 30079
rect 356 30045 430 30079
rect 245 30011 430 30045
rect 245 29977 322 30011
rect 356 29977 430 30011
rect 245 29943 430 29977
rect 245 29909 322 29943
rect 356 29909 430 29943
rect 245 29875 430 29909
rect 245 29841 322 29875
rect 356 29841 430 29875
rect 245 29807 430 29841
rect 245 29773 322 29807
rect 356 29773 430 29807
rect 245 29739 430 29773
rect 245 29705 322 29739
rect 356 29705 430 29739
rect 245 29671 430 29705
rect 245 29637 322 29671
rect 356 29637 430 29671
rect 245 29603 430 29637
rect 245 29569 322 29603
rect 356 29569 430 29603
rect 245 29535 430 29569
rect 245 29501 322 29535
rect 356 29501 430 29535
rect 245 29467 430 29501
rect 245 29433 322 29467
rect 356 29433 430 29467
rect 245 29399 430 29433
rect 245 29365 322 29399
rect 356 29365 430 29399
rect 245 29331 430 29365
rect 245 29297 322 29331
rect 356 29297 430 29331
rect 245 29263 430 29297
rect 245 29229 322 29263
rect 356 29229 430 29263
rect 245 29195 430 29229
rect 245 29161 322 29195
rect 356 29161 430 29195
rect 245 29127 430 29161
rect 245 29093 322 29127
rect 356 29093 430 29127
rect 245 29059 430 29093
rect 245 29025 322 29059
rect 356 29025 430 29059
rect 245 28991 430 29025
rect 245 28957 322 28991
rect 356 28957 430 28991
rect 245 28923 430 28957
rect 245 28889 322 28923
rect 356 28889 430 28923
rect 245 28855 430 28889
rect 245 28821 322 28855
rect 356 28821 430 28855
rect 245 28787 430 28821
rect 245 28753 322 28787
rect 356 28753 430 28787
rect 245 28719 430 28753
rect 245 28685 322 28719
rect 356 28685 430 28719
rect 245 28651 430 28685
rect 245 28617 322 28651
rect 356 28617 430 28651
rect 245 28583 430 28617
rect 245 28549 322 28583
rect 356 28549 430 28583
rect 245 28515 430 28549
rect 245 28481 322 28515
rect 356 28481 430 28515
rect 245 28447 430 28481
rect 245 28413 322 28447
rect 356 28413 430 28447
rect 245 28379 430 28413
rect 245 28345 322 28379
rect 356 28345 430 28379
rect 245 28311 430 28345
rect 245 28277 322 28311
rect 356 28277 430 28311
rect 245 28243 430 28277
rect 245 28209 322 28243
rect 356 28209 430 28243
rect 245 28175 430 28209
rect 245 28141 322 28175
rect 356 28141 430 28175
rect 245 28107 430 28141
rect 245 28073 322 28107
rect 356 28073 430 28107
rect 245 28039 430 28073
rect 245 28005 322 28039
rect 356 28005 430 28039
rect 245 27971 430 28005
rect 245 27937 322 27971
rect 356 27937 430 27971
rect 245 27903 430 27937
rect 245 27869 322 27903
rect 356 27869 430 27903
rect 245 27835 430 27869
rect 245 27801 322 27835
rect 356 27801 430 27835
rect 245 27767 430 27801
rect 245 27733 322 27767
rect 356 27733 430 27767
rect 245 27699 430 27733
rect 245 27665 322 27699
rect 356 27665 430 27699
rect 245 27631 430 27665
rect 245 27597 322 27631
rect 356 27597 430 27631
rect 245 27563 430 27597
rect 245 27529 322 27563
rect 356 27529 430 27563
rect 245 27495 430 27529
rect 245 27461 322 27495
rect 356 27461 430 27495
rect 245 27427 430 27461
rect 245 27393 322 27427
rect 356 27393 430 27427
rect 245 27359 430 27393
rect 245 27325 322 27359
rect 356 27325 430 27359
rect 245 27291 430 27325
rect 245 27257 322 27291
rect 356 27257 430 27291
rect 245 27223 430 27257
rect 245 27189 322 27223
rect 356 27189 430 27223
rect 245 27155 430 27189
rect 245 27121 322 27155
rect 356 27121 430 27155
rect 245 27087 430 27121
rect 245 27053 322 27087
rect 356 27053 430 27087
rect 245 27019 430 27053
rect 245 26985 322 27019
rect 356 26985 430 27019
rect 245 26951 430 26985
rect 245 26917 322 26951
rect 356 26917 430 26951
rect 245 26883 430 26917
rect 245 26849 322 26883
rect 356 26849 430 26883
rect 245 26815 430 26849
rect 245 26781 322 26815
rect 356 26781 430 26815
rect 245 26747 430 26781
rect 245 26713 322 26747
rect 356 26713 430 26747
rect 245 26679 430 26713
rect 245 26645 322 26679
rect 356 26645 430 26679
rect 245 26611 430 26645
rect 245 26577 322 26611
rect 356 26577 430 26611
rect 245 26543 430 26577
rect 245 26509 322 26543
rect 356 26509 430 26543
rect 245 26475 430 26509
rect 245 26441 322 26475
rect 356 26441 430 26475
rect 245 26407 430 26441
rect 245 26373 322 26407
rect 356 26373 430 26407
rect 245 26339 430 26373
rect 245 26305 322 26339
rect 356 26305 430 26339
rect 245 26271 430 26305
rect 245 26237 322 26271
rect 356 26237 430 26271
rect 245 26203 430 26237
rect 245 26169 322 26203
rect 356 26169 430 26203
rect 245 26135 430 26169
rect 245 26101 322 26135
rect 356 26101 430 26135
rect 245 26067 430 26101
rect 245 26033 322 26067
rect 356 26033 430 26067
rect 245 25999 430 26033
rect 245 25965 322 25999
rect 356 25965 430 25999
rect 245 25931 430 25965
rect 245 25897 322 25931
rect 356 25897 430 25931
rect 245 25863 430 25897
rect 245 25829 322 25863
rect 356 25829 430 25863
rect 245 25795 430 25829
rect 245 25761 322 25795
rect 356 25761 430 25795
rect 245 25727 430 25761
rect 245 25693 322 25727
rect 356 25693 430 25727
rect 245 25659 430 25693
rect 245 25625 322 25659
rect 356 25625 430 25659
rect 245 25591 430 25625
rect 245 25557 322 25591
rect 356 25557 430 25591
rect 245 25523 430 25557
rect 245 25489 322 25523
rect 356 25489 430 25523
rect 245 25455 430 25489
rect 245 25421 322 25455
rect 356 25421 430 25455
rect 245 25387 430 25421
rect 245 25353 322 25387
rect 356 25353 430 25387
rect 245 25319 430 25353
rect 245 25285 322 25319
rect 356 25285 430 25319
rect 245 25251 430 25285
rect 245 25217 322 25251
rect 356 25217 430 25251
rect 245 25183 430 25217
rect 245 25149 322 25183
rect 356 25149 430 25183
rect 245 25115 430 25149
rect 245 25081 322 25115
rect 356 25081 430 25115
rect 245 25047 430 25081
rect 245 25013 322 25047
rect 356 25013 430 25047
rect 245 24979 430 25013
rect 245 24945 322 24979
rect 356 24945 430 24979
rect 245 24911 430 24945
rect 245 24877 322 24911
rect 356 24877 430 24911
rect 245 24843 430 24877
rect 245 24809 322 24843
rect 356 24809 430 24843
rect 245 24775 430 24809
rect 245 24741 322 24775
rect 356 24741 430 24775
rect 245 24707 430 24741
rect 245 24673 322 24707
rect 356 24673 430 24707
rect 245 24639 430 24673
rect 245 24605 322 24639
rect 356 24605 430 24639
rect 245 24571 430 24605
rect 245 24537 322 24571
rect 356 24537 430 24571
rect 245 24503 430 24537
rect 245 24469 322 24503
rect 356 24469 430 24503
rect 245 24435 430 24469
rect 245 24401 322 24435
rect 356 24401 430 24435
rect 245 24367 430 24401
rect 245 24333 322 24367
rect 356 24333 430 24367
rect 245 24299 430 24333
rect 245 24265 322 24299
rect 356 24265 430 24299
rect 245 24231 430 24265
rect 245 24197 322 24231
rect 356 24197 430 24231
rect 245 24163 430 24197
rect 245 24129 322 24163
rect 356 24129 430 24163
rect 245 24095 430 24129
rect 245 24061 322 24095
rect 356 24061 430 24095
rect 245 24027 430 24061
rect 245 23993 322 24027
rect 356 23993 430 24027
rect 245 23959 430 23993
rect 245 23925 322 23959
rect 356 23925 430 23959
rect 245 23891 430 23925
rect 245 23857 322 23891
rect 356 23857 430 23891
rect 245 23823 430 23857
rect 245 23789 322 23823
rect 356 23789 430 23823
rect 245 23755 430 23789
rect 245 23721 322 23755
rect 356 23721 430 23755
rect 245 23687 430 23721
rect 245 23653 322 23687
rect 356 23653 430 23687
rect 245 23619 430 23653
rect 245 23585 322 23619
rect 356 23585 430 23619
rect 245 23551 430 23585
rect 245 23517 322 23551
rect 356 23517 430 23551
rect 245 23483 430 23517
rect 245 23449 322 23483
rect 356 23449 430 23483
rect 245 23415 430 23449
rect 245 23381 322 23415
rect 356 23381 430 23415
rect 245 23347 430 23381
rect 245 23313 322 23347
rect 356 23313 430 23347
rect 245 23279 430 23313
rect 245 23245 322 23279
rect 356 23245 430 23279
rect 245 23211 430 23245
rect 245 23177 322 23211
rect 356 23177 430 23211
rect 245 23143 430 23177
rect 245 23109 322 23143
rect 356 23109 430 23143
rect 245 23075 430 23109
rect 245 23041 322 23075
rect 356 23041 430 23075
rect 245 23007 430 23041
rect 245 22973 322 23007
rect 356 22973 430 23007
rect 245 22939 430 22973
rect 245 22905 322 22939
rect 356 22905 430 22939
rect 245 22871 430 22905
rect 245 22837 322 22871
rect 356 22837 430 22871
rect 245 22803 430 22837
rect 245 22769 322 22803
rect 356 22769 430 22803
rect 245 22735 430 22769
rect 245 22701 322 22735
rect 356 22701 430 22735
rect 245 22667 430 22701
rect 245 22633 322 22667
rect 356 22633 430 22667
rect 245 22599 430 22633
rect 245 22565 322 22599
rect 356 22565 430 22599
rect 245 22531 430 22565
rect 245 22497 322 22531
rect 356 22497 430 22531
rect 245 22463 430 22497
rect 245 22429 322 22463
rect 356 22429 430 22463
rect 245 22395 430 22429
rect 245 22361 322 22395
rect 356 22361 430 22395
rect 245 22327 430 22361
rect 245 22293 322 22327
rect 356 22293 430 22327
rect 245 22259 430 22293
rect 245 22225 322 22259
rect 356 22225 430 22259
rect 245 22191 430 22225
rect 245 22157 322 22191
rect 356 22157 430 22191
rect 245 22123 430 22157
rect 245 22089 322 22123
rect 356 22089 430 22123
rect 245 22055 430 22089
rect 245 22021 322 22055
rect 356 22021 430 22055
rect 245 21987 430 22021
rect 245 21953 322 21987
rect 356 21953 430 21987
rect 245 21919 430 21953
rect 245 21885 322 21919
rect 356 21885 430 21919
rect 245 21851 430 21885
rect 245 21817 322 21851
rect 356 21817 430 21851
rect 245 21783 430 21817
rect 245 21749 322 21783
rect 356 21749 430 21783
rect 245 21715 430 21749
rect 245 21681 322 21715
rect 356 21681 430 21715
rect 245 21647 430 21681
rect 245 21613 322 21647
rect 356 21613 430 21647
rect 245 21579 430 21613
rect 245 21545 322 21579
rect 356 21545 430 21579
rect 245 21511 430 21545
rect 245 21477 322 21511
rect 356 21477 430 21511
rect 245 21443 430 21477
rect 245 21409 322 21443
rect 356 21409 430 21443
rect 245 21375 430 21409
rect 245 21341 322 21375
rect 356 21341 430 21375
rect 245 21307 430 21341
rect 245 21273 322 21307
rect 356 21273 430 21307
rect 245 21239 430 21273
rect 245 21205 322 21239
rect 356 21205 430 21239
rect 245 21171 430 21205
rect 245 21137 322 21171
rect 356 21137 430 21171
rect 245 21103 430 21137
rect 245 21069 322 21103
rect 356 21069 430 21103
rect 245 21035 430 21069
rect 245 21001 322 21035
rect 356 21001 430 21035
rect 245 20967 430 21001
rect 245 20933 322 20967
rect 356 20933 430 20967
rect 245 20899 430 20933
rect 245 20865 322 20899
rect 356 20865 430 20899
rect 245 20831 430 20865
rect 245 20797 322 20831
rect 356 20797 430 20831
rect 245 20763 430 20797
rect 245 20729 322 20763
rect 356 20729 430 20763
rect 245 20695 430 20729
rect 245 20661 322 20695
rect 356 20661 430 20695
rect 245 20627 430 20661
rect 245 20593 322 20627
rect 356 20593 430 20627
rect 245 20559 430 20593
rect 245 20525 322 20559
rect 356 20525 430 20559
rect 245 20491 430 20525
rect 245 20457 322 20491
rect 356 20457 430 20491
rect 245 20423 430 20457
rect 245 20389 322 20423
rect 356 20389 430 20423
rect 245 20355 430 20389
rect 245 20321 322 20355
rect 356 20321 430 20355
rect 245 20287 430 20321
rect 245 20253 322 20287
rect 356 20253 430 20287
rect 245 20219 430 20253
rect 245 20185 322 20219
rect 356 20185 430 20219
rect 245 20151 430 20185
rect 245 20117 322 20151
rect 356 20117 430 20151
rect 245 20083 430 20117
rect 245 20049 322 20083
rect 356 20049 430 20083
rect 245 20015 430 20049
rect 245 19981 322 20015
rect 356 19981 430 20015
rect 245 19947 430 19981
rect 245 19913 322 19947
rect 356 19913 430 19947
rect 245 19879 430 19913
rect 245 19845 322 19879
rect 356 19845 430 19879
rect 245 19811 430 19845
rect 245 19777 322 19811
rect 356 19777 430 19811
rect 245 19743 430 19777
rect 245 19709 322 19743
rect 356 19709 430 19743
rect 245 19675 430 19709
rect 245 19641 322 19675
rect 356 19641 430 19675
rect 245 19607 430 19641
rect 245 19573 322 19607
rect 356 19573 430 19607
rect 245 19539 430 19573
rect 245 19505 322 19539
rect 356 19505 430 19539
rect 245 19471 430 19505
rect 245 19437 322 19471
rect 356 19437 430 19471
rect 245 19403 430 19437
rect 245 19369 322 19403
rect 356 19369 430 19403
rect 245 19335 430 19369
rect 245 19301 322 19335
rect 356 19301 430 19335
rect 245 19267 430 19301
rect 245 19233 322 19267
rect 356 19233 430 19267
rect 245 19199 430 19233
rect 245 19165 322 19199
rect 356 19165 430 19199
rect 245 19131 430 19165
rect 245 19097 322 19131
rect 356 19097 430 19131
rect 245 19063 430 19097
rect 245 19029 322 19063
rect 356 19029 430 19063
rect 245 18995 430 19029
rect 245 18961 322 18995
rect 356 18961 430 18995
rect 245 18927 430 18961
rect 245 18893 322 18927
rect 356 18893 430 18927
rect 245 18859 430 18893
rect 245 18825 322 18859
rect 356 18825 430 18859
rect 245 18791 430 18825
rect 245 18757 322 18791
rect 356 18757 430 18791
rect 245 18723 430 18757
rect 245 18689 322 18723
rect 356 18689 430 18723
rect 245 18655 430 18689
rect 245 18621 322 18655
rect 356 18621 430 18655
rect 245 18587 430 18621
rect 245 18553 322 18587
rect 356 18553 430 18587
rect 245 18519 430 18553
rect 245 18485 322 18519
rect 356 18485 430 18519
rect 245 18451 430 18485
rect 245 18417 322 18451
rect 356 18417 430 18451
rect 245 18383 430 18417
rect 245 18349 322 18383
rect 356 18349 430 18383
rect 245 18315 430 18349
rect 245 18281 322 18315
rect 356 18281 430 18315
rect 245 18247 430 18281
rect 245 18213 322 18247
rect 356 18213 430 18247
rect 245 18179 430 18213
rect 245 18145 322 18179
rect 356 18145 430 18179
rect 245 18111 430 18145
rect 245 18077 322 18111
rect 356 18077 430 18111
rect 245 18043 430 18077
rect 245 18009 322 18043
rect 356 18009 430 18043
rect 245 17975 430 18009
rect 245 17941 322 17975
rect 356 17941 430 17975
rect 245 17907 430 17941
rect 245 17873 322 17907
rect 356 17873 430 17907
rect 245 17839 430 17873
rect 245 17805 322 17839
rect 356 17805 430 17839
rect 245 17771 430 17805
rect 245 17737 322 17771
rect 356 17737 430 17771
rect 245 17703 430 17737
rect 245 17669 322 17703
rect 356 17669 430 17703
rect 245 17635 430 17669
rect 245 17601 322 17635
rect 356 17601 430 17635
rect 245 17567 430 17601
rect 245 17533 322 17567
rect 356 17533 430 17567
rect 245 17499 430 17533
rect 245 17465 322 17499
rect 356 17465 430 17499
rect 245 17431 430 17465
rect 245 17397 322 17431
rect 356 17397 430 17431
rect 245 17363 430 17397
rect 245 17329 322 17363
rect 356 17329 430 17363
rect 245 17295 430 17329
rect 245 17261 322 17295
rect 356 17261 430 17295
rect 245 17227 430 17261
rect 245 17193 322 17227
rect 356 17193 430 17227
rect 245 17159 430 17193
rect 245 17125 322 17159
rect 356 17125 430 17159
rect 245 17091 430 17125
rect 245 17057 322 17091
rect 356 17057 430 17091
rect 245 17023 430 17057
rect 245 16989 322 17023
rect 356 16989 430 17023
rect 245 16955 430 16989
rect 245 16921 322 16955
rect 356 16921 430 16955
rect 245 16887 430 16921
rect 245 16853 322 16887
rect 356 16853 430 16887
rect 245 16819 430 16853
rect 245 16785 322 16819
rect 356 16785 430 16819
rect 245 16751 430 16785
rect 245 16717 322 16751
rect 356 16717 430 16751
rect 245 16683 430 16717
rect 245 16649 322 16683
rect 356 16649 430 16683
rect 245 16615 430 16649
rect 245 16581 322 16615
rect 356 16581 430 16615
rect 245 16547 430 16581
rect 245 16513 322 16547
rect 356 16513 430 16547
rect 245 16479 430 16513
rect 245 16445 322 16479
rect 356 16445 430 16479
rect 245 16411 430 16445
rect 245 16377 322 16411
rect 356 16377 430 16411
rect 245 16343 430 16377
rect 245 16309 322 16343
rect 356 16309 430 16343
rect 245 16275 430 16309
rect 245 16241 322 16275
rect 356 16241 430 16275
rect 245 16207 430 16241
rect 245 16173 322 16207
rect 356 16173 430 16207
rect 245 16139 430 16173
rect 245 16105 322 16139
rect 356 16105 430 16139
rect 245 16071 430 16105
rect 245 16037 322 16071
rect 356 16037 430 16071
rect 245 16003 430 16037
rect 245 15969 322 16003
rect 356 15969 430 16003
rect 245 15935 430 15969
rect 245 15901 322 15935
rect 356 15901 430 15935
rect 245 15867 430 15901
rect 245 15833 322 15867
rect 356 15833 430 15867
rect 245 15799 430 15833
rect 245 15765 322 15799
rect 356 15765 430 15799
rect 245 15731 430 15765
rect 245 15697 322 15731
rect 356 15697 430 15731
rect 245 15663 430 15697
rect 245 15629 322 15663
rect 356 15629 430 15663
rect 245 15595 430 15629
rect 245 15561 322 15595
rect 356 15561 430 15595
rect 245 15527 430 15561
rect 245 15493 322 15527
rect 356 15493 430 15527
rect 245 15459 430 15493
rect 245 15425 322 15459
rect 356 15425 430 15459
rect 245 15391 430 15425
rect 245 15357 322 15391
rect 356 15357 430 15391
rect 245 15323 430 15357
rect 245 15289 322 15323
rect 356 15289 430 15323
rect 245 15255 430 15289
rect 245 15221 322 15255
rect 356 15221 430 15255
rect 245 15187 430 15221
rect 245 15153 322 15187
rect 356 15153 430 15187
rect 245 15119 430 15153
rect 245 15085 322 15119
rect 356 15085 430 15119
rect 245 15051 430 15085
rect 245 15017 322 15051
rect 356 15017 430 15051
rect 245 14983 430 15017
rect 245 14949 322 14983
rect 356 14949 430 14983
rect 245 14915 430 14949
rect 245 14881 322 14915
rect 356 14881 430 14915
rect 245 14847 430 14881
rect 245 14813 322 14847
rect 356 14813 430 14847
rect 245 14779 430 14813
rect 245 14745 322 14779
rect 356 14745 430 14779
rect 245 14711 430 14745
rect 245 14677 322 14711
rect 356 14677 430 14711
rect 245 14643 430 14677
rect 245 14609 322 14643
rect 356 14609 430 14643
rect 245 14575 430 14609
rect 245 14541 322 14575
rect 356 14541 430 14575
rect 245 14507 430 14541
rect 245 14473 322 14507
rect 356 14473 430 14507
rect 245 14439 430 14473
rect 245 14405 322 14439
rect 356 14405 430 14439
rect 245 14371 430 14405
rect 245 14337 322 14371
rect 356 14337 430 14371
rect 245 14303 430 14337
rect 245 14269 322 14303
rect 356 14269 430 14303
rect 245 14235 430 14269
rect 245 14201 322 14235
rect 356 14201 430 14235
rect 245 14167 430 14201
rect 245 14133 322 14167
rect 356 14133 430 14167
rect 245 14099 430 14133
rect 245 14065 322 14099
rect 356 14065 430 14099
rect 245 14031 430 14065
rect 245 13997 322 14031
rect 356 13997 430 14031
rect 245 13963 430 13997
rect 245 13929 322 13963
rect 356 13929 430 13963
rect 245 13895 430 13929
rect 245 13861 322 13895
rect 356 13861 430 13895
rect 245 13827 430 13861
rect 245 13793 322 13827
rect 356 13793 430 13827
rect 245 13759 430 13793
rect 245 13725 322 13759
rect 356 13725 430 13759
rect 245 13691 430 13725
rect 245 13657 322 13691
rect 356 13657 430 13691
rect 245 13623 430 13657
rect 245 13589 322 13623
rect 356 13589 430 13623
rect 245 13555 430 13589
rect 245 13521 322 13555
rect 356 13521 430 13555
rect 245 13487 430 13521
rect 245 13453 322 13487
rect 356 13453 430 13487
rect 245 13419 430 13453
rect 245 13385 322 13419
rect 356 13385 430 13419
rect 245 13351 430 13385
rect 245 13317 322 13351
rect 356 13317 430 13351
rect 245 13283 430 13317
rect 245 13249 322 13283
rect 356 13249 430 13283
rect 245 13215 430 13249
rect 245 13181 322 13215
rect 356 13181 430 13215
rect 245 13147 430 13181
rect 245 13113 322 13147
rect 356 13113 430 13147
rect 245 13079 430 13113
rect 245 13045 322 13079
rect 356 13045 430 13079
rect 245 13011 430 13045
rect 245 12977 322 13011
rect 356 12977 430 13011
rect 245 12943 430 12977
rect 245 12909 322 12943
rect 356 12909 430 12943
rect 245 12875 430 12909
rect 245 12841 322 12875
rect 356 12841 430 12875
rect 245 12807 430 12841
rect 245 12773 322 12807
rect 356 12773 430 12807
rect 245 12739 430 12773
rect 245 12705 322 12739
rect 356 12705 430 12739
rect 245 12671 430 12705
rect 245 12637 322 12671
rect 356 12637 430 12671
rect 245 12603 430 12637
rect 245 12569 322 12603
rect 356 12569 430 12603
rect 245 12535 430 12569
rect 245 12501 322 12535
rect 356 12501 430 12535
rect 245 12467 430 12501
rect 245 12433 322 12467
rect 356 12433 430 12467
rect 245 12399 430 12433
rect 245 12365 322 12399
rect 356 12365 430 12399
rect 245 12331 430 12365
rect 245 12297 322 12331
rect 356 12297 430 12331
rect 245 12263 430 12297
rect 245 12229 322 12263
rect 356 12229 430 12263
rect 245 12195 430 12229
rect 245 12161 322 12195
rect 356 12161 430 12195
rect 245 12127 430 12161
rect 245 12093 322 12127
rect 356 12093 430 12127
rect 245 12059 430 12093
rect 245 12025 322 12059
rect 356 12025 430 12059
rect 245 11991 430 12025
rect 245 11957 322 11991
rect 356 11957 430 11991
rect 245 11923 430 11957
rect 245 11889 322 11923
rect 356 11889 430 11923
rect 245 11855 430 11889
rect 245 11821 322 11855
rect 356 11821 430 11855
rect 245 11787 430 11821
rect 245 11753 322 11787
rect 356 11753 430 11787
rect 245 11719 430 11753
rect 245 11685 322 11719
rect 356 11685 430 11719
rect 245 11651 430 11685
rect 245 11617 322 11651
rect 356 11617 430 11651
rect 245 11583 430 11617
rect 245 11549 322 11583
rect 356 11549 430 11583
rect 245 11515 430 11549
rect 245 11481 322 11515
rect 356 11481 430 11515
rect 245 11447 430 11481
rect 245 11413 322 11447
rect 356 11413 430 11447
rect 245 11379 430 11413
rect 245 11345 322 11379
rect 356 11345 430 11379
rect 245 11311 430 11345
rect 245 11277 322 11311
rect 356 11277 430 11311
rect 245 11243 430 11277
rect 245 11209 322 11243
rect 356 11209 430 11243
rect 245 11175 430 11209
rect 245 11141 322 11175
rect 356 11141 430 11175
rect 245 11107 430 11141
rect 245 11073 322 11107
rect 356 11073 430 11107
rect 245 11039 430 11073
rect 245 11005 322 11039
rect 356 11005 430 11039
rect 245 10971 430 11005
rect 245 10937 322 10971
rect 356 10937 430 10971
rect 245 10903 430 10937
rect 245 10869 322 10903
rect 356 10869 430 10903
rect 245 10835 430 10869
rect 245 10801 322 10835
rect 356 10801 430 10835
rect 245 10767 430 10801
rect 245 10733 322 10767
rect 356 10733 430 10767
rect 245 10699 430 10733
rect 245 10665 322 10699
rect 356 10665 430 10699
rect 245 10631 430 10665
rect 245 10597 322 10631
rect 356 10597 430 10631
rect 245 10563 430 10597
rect 245 10529 322 10563
rect 356 10529 430 10563
rect 245 10495 430 10529
rect 245 10461 322 10495
rect 356 10461 430 10495
rect 245 10427 430 10461
rect 245 10393 322 10427
rect 356 10393 430 10427
rect 245 10359 430 10393
rect 245 10325 322 10359
rect 356 10325 430 10359
rect 245 10291 430 10325
rect 245 10257 322 10291
rect 356 10257 430 10291
rect 245 10223 430 10257
rect 245 10189 322 10223
rect 356 10189 430 10223
rect 245 10155 430 10189
rect 245 10121 322 10155
rect 356 10121 430 10155
rect 245 10087 430 10121
rect 245 10053 322 10087
rect 356 10053 430 10087
rect 245 10019 430 10053
rect 245 9985 322 10019
rect 356 9985 430 10019
rect 245 9951 430 9985
rect 245 9917 322 9951
rect 356 9917 430 9951
rect 245 9883 430 9917
rect 245 9849 322 9883
rect 356 9849 430 9883
rect 245 9815 430 9849
rect 245 9781 322 9815
rect 356 9781 430 9815
rect 245 9747 430 9781
rect 245 9713 322 9747
rect 356 9713 430 9747
rect 245 9679 430 9713
rect 1177 34636 13817 34684
rect 1177 34602 1365 34636
rect 1399 34602 1433 34636
rect 1467 34602 1501 34636
rect 1535 34602 1569 34636
rect 1603 34602 1637 34636
rect 1671 34602 1705 34636
rect 1739 34602 1773 34636
rect 1807 34602 1841 34636
rect 1875 34602 1909 34636
rect 1943 34602 1977 34636
rect 2011 34602 2045 34636
rect 2079 34602 2113 34636
rect 2147 34602 2181 34636
rect 2215 34602 2249 34636
rect 2283 34602 2317 34636
rect 2351 34602 2385 34636
rect 2419 34602 2453 34636
rect 2487 34602 2521 34636
rect 2555 34602 2589 34636
rect 2623 34602 2657 34636
rect 2691 34602 2725 34636
rect 2759 34602 2793 34636
rect 2827 34602 2861 34636
rect 2895 34602 2929 34636
rect 2963 34602 2997 34636
rect 3031 34602 3065 34636
rect 3099 34602 3133 34636
rect 3167 34602 3201 34636
rect 3235 34602 3269 34636
rect 3303 34602 3337 34636
rect 3371 34602 3405 34636
rect 3439 34602 3473 34636
rect 3507 34602 3541 34636
rect 3575 34602 3609 34636
rect 3643 34602 3677 34636
rect 3711 34602 3745 34636
rect 3779 34602 3813 34636
rect 3847 34602 3881 34636
rect 3915 34602 3949 34636
rect 3983 34602 4017 34636
rect 4051 34602 4085 34636
rect 4119 34602 4153 34636
rect 4187 34602 4221 34636
rect 4255 34602 4289 34636
rect 4323 34602 4357 34636
rect 4391 34602 4425 34636
rect 4459 34602 4493 34636
rect 4527 34602 4561 34636
rect 4595 34602 4629 34636
rect 4663 34602 4697 34636
rect 4731 34602 4765 34636
rect 4799 34602 4833 34636
rect 4867 34602 4901 34636
rect 4935 34602 4969 34636
rect 5003 34602 5037 34636
rect 5071 34602 5105 34636
rect 5139 34602 5173 34636
rect 5207 34602 5241 34636
rect 5275 34602 5309 34636
rect 5343 34602 5377 34636
rect 5411 34602 5445 34636
rect 5479 34602 5513 34636
rect 5547 34602 5581 34636
rect 5615 34602 5649 34636
rect 5683 34602 5717 34636
rect 5751 34602 5785 34636
rect 5819 34602 5853 34636
rect 5887 34602 5921 34636
rect 5955 34602 5989 34636
rect 6023 34602 6057 34636
rect 6091 34602 6125 34636
rect 6159 34602 6193 34636
rect 6227 34602 6261 34636
rect 6295 34602 6329 34636
rect 6363 34602 6397 34636
rect 6431 34602 6465 34636
rect 6499 34602 6533 34636
rect 6567 34602 6601 34636
rect 6635 34602 6669 34636
rect 6703 34602 6737 34636
rect 6771 34602 6805 34636
rect 6839 34602 6873 34636
rect 6907 34602 6941 34636
rect 6975 34602 7009 34636
rect 7043 34602 7077 34636
rect 7111 34602 7145 34636
rect 7179 34602 7213 34636
rect 7247 34602 7281 34636
rect 7315 34602 7349 34636
rect 7383 34602 7417 34636
rect 7451 34602 7485 34636
rect 7519 34602 7553 34636
rect 7587 34602 7621 34636
rect 7655 34602 7689 34636
rect 7723 34602 7757 34636
rect 7791 34602 7825 34636
rect 7859 34602 7893 34636
rect 7927 34602 7961 34636
rect 7995 34602 8029 34636
rect 8063 34602 8097 34636
rect 8131 34602 8165 34636
rect 8199 34602 8233 34636
rect 8267 34602 8301 34636
rect 8335 34602 8369 34636
rect 8403 34602 8437 34636
rect 8471 34602 8505 34636
rect 8539 34602 8573 34636
rect 8607 34602 8641 34636
rect 8675 34602 8709 34636
rect 8743 34602 8777 34636
rect 8811 34602 8845 34636
rect 8879 34602 8913 34636
rect 8947 34602 8981 34636
rect 9015 34602 9049 34636
rect 9083 34602 9117 34636
rect 9151 34602 9185 34636
rect 9219 34602 9253 34636
rect 9287 34602 9321 34636
rect 9355 34602 9389 34636
rect 9423 34602 9457 34636
rect 9491 34602 9525 34636
rect 9559 34602 9593 34636
rect 9627 34602 9661 34636
rect 9695 34602 9729 34636
rect 9763 34602 9797 34636
rect 9831 34602 9865 34636
rect 9899 34602 9933 34636
rect 9967 34602 10001 34636
rect 10035 34602 10069 34636
rect 10103 34602 10137 34636
rect 10171 34602 10205 34636
rect 10239 34602 10273 34636
rect 10307 34602 10341 34636
rect 10375 34602 10409 34636
rect 10443 34602 10477 34636
rect 10511 34602 10545 34636
rect 10579 34602 10613 34636
rect 10647 34602 10681 34636
rect 10715 34602 10749 34636
rect 10783 34602 10817 34636
rect 10851 34602 10885 34636
rect 10919 34602 10953 34636
rect 10987 34602 11021 34636
rect 11055 34602 11089 34636
rect 11123 34602 11157 34636
rect 11191 34602 11225 34636
rect 11259 34602 11293 34636
rect 11327 34602 11361 34636
rect 11395 34602 11429 34636
rect 11463 34602 11497 34636
rect 11531 34602 11565 34636
rect 11599 34602 11633 34636
rect 11667 34602 11701 34636
rect 11735 34602 11769 34636
rect 11803 34602 11837 34636
rect 11871 34602 11905 34636
rect 11939 34602 11973 34636
rect 12007 34602 12041 34636
rect 12075 34602 12109 34636
rect 12143 34602 12177 34636
rect 12211 34602 12245 34636
rect 12279 34602 12313 34636
rect 12347 34602 12381 34636
rect 12415 34602 12449 34636
rect 12483 34602 12517 34636
rect 12551 34602 12585 34636
rect 12619 34602 12653 34636
rect 12687 34602 12721 34636
rect 12755 34602 12789 34636
rect 12823 34602 12857 34636
rect 12891 34602 12925 34636
rect 12959 34602 12993 34636
rect 13027 34602 13061 34636
rect 13095 34602 13129 34636
rect 13163 34602 13197 34636
rect 13231 34602 13265 34636
rect 13299 34602 13333 34636
rect 13367 34602 13401 34636
rect 13435 34602 13469 34636
rect 13503 34602 13537 34636
rect 13571 34602 13605 34636
rect 13639 34602 13817 34636
rect 1177 34564 13817 34602
rect 1177 34486 1297 34564
rect 1177 34452 1221 34486
rect 1255 34452 1297 34486
rect 1177 34418 1297 34452
rect 1177 34384 1221 34418
rect 1255 34384 1297 34418
rect 1177 34350 1297 34384
rect 1177 34316 1221 34350
rect 1255 34316 1297 34350
rect 1177 34282 1297 34316
rect 1177 34248 1221 34282
rect 1255 34248 1297 34282
rect 1177 34214 1297 34248
rect 1177 34180 1221 34214
rect 1255 34180 1297 34214
rect 1177 34146 1297 34180
rect 1177 34112 1221 34146
rect 1255 34112 1297 34146
rect 1177 34078 1297 34112
rect 1177 34044 1221 34078
rect 1255 34044 1297 34078
rect 1177 34010 1297 34044
rect 1177 33976 1221 34010
rect 1255 33976 1297 34010
rect 1177 33942 1297 33976
rect 1177 33908 1221 33942
rect 1255 33908 1297 33942
rect 1177 33874 1297 33908
rect 1177 33840 1221 33874
rect 1255 33840 1297 33874
rect 1177 33806 1297 33840
rect 1177 33772 1221 33806
rect 1255 33772 1297 33806
rect 1177 33738 1297 33772
rect 1177 33704 1221 33738
rect 1255 33704 1297 33738
rect 1177 33670 1297 33704
rect 1177 33636 1221 33670
rect 1255 33636 1297 33670
rect 1177 33602 1297 33636
rect 1177 33568 1221 33602
rect 1255 33568 1297 33602
rect 1177 33534 1297 33568
rect 1177 33500 1221 33534
rect 1255 33500 1297 33534
rect 1177 33466 1297 33500
rect 1177 33432 1221 33466
rect 1255 33432 1297 33466
rect 1177 33398 1297 33432
rect 1177 33364 1221 33398
rect 1255 33364 1297 33398
rect 1177 33330 1297 33364
rect 1177 33296 1221 33330
rect 1255 33296 1297 33330
rect 1177 33262 1297 33296
rect 1177 33228 1221 33262
rect 1255 33228 1297 33262
rect 1177 33194 1297 33228
rect 1177 33160 1221 33194
rect 1255 33160 1297 33194
rect 1177 33126 1297 33160
rect 1177 33092 1221 33126
rect 1255 33092 1297 33126
rect 1177 33058 1297 33092
rect 1177 33024 1221 33058
rect 1255 33024 1297 33058
rect 1177 32990 1297 33024
rect 1177 32956 1221 32990
rect 1255 32956 1297 32990
rect 1177 32922 1297 32956
rect 1177 32888 1221 32922
rect 1255 32888 1297 32922
rect 1177 32854 1297 32888
rect 1177 32820 1221 32854
rect 1255 32820 1297 32854
rect 1177 32786 1297 32820
rect 1177 32752 1221 32786
rect 1255 32752 1297 32786
rect 1177 32718 1297 32752
rect 1177 32684 1221 32718
rect 1255 32684 1297 32718
rect 1177 32650 1297 32684
rect 1177 32616 1221 32650
rect 1255 32616 1297 32650
rect 1177 32582 1297 32616
rect 1177 32548 1221 32582
rect 1255 32548 1297 32582
rect 1177 32514 1297 32548
rect 1177 32480 1221 32514
rect 1255 32480 1297 32514
rect 1177 32446 1297 32480
rect 1177 32412 1221 32446
rect 1255 32412 1297 32446
rect 1177 32378 1297 32412
rect 1177 32344 1221 32378
rect 1255 32344 1297 32378
rect 1177 32310 1297 32344
rect 1177 32276 1221 32310
rect 1255 32276 1297 32310
rect 1177 32242 1297 32276
rect 1177 32208 1221 32242
rect 1255 32208 1297 32242
rect 1177 32174 1297 32208
rect 1177 32140 1221 32174
rect 1255 32140 1297 32174
rect 1177 32106 1297 32140
rect 1177 32072 1221 32106
rect 1255 32072 1297 32106
rect 1177 32038 1297 32072
rect 1177 32004 1221 32038
rect 1255 32004 1297 32038
rect 1177 31970 1297 32004
rect 1177 31936 1221 31970
rect 1255 31936 1297 31970
rect 1177 31902 1297 31936
rect 1177 31868 1221 31902
rect 1255 31868 1297 31902
rect 1177 31834 1297 31868
rect 1177 31800 1221 31834
rect 1255 31800 1297 31834
rect 1177 31766 1297 31800
rect 1177 31732 1221 31766
rect 1255 31732 1297 31766
rect 1177 31698 1297 31732
rect 1177 31664 1221 31698
rect 1255 31664 1297 31698
rect 1177 31630 1297 31664
rect 1177 31596 1221 31630
rect 1255 31596 1297 31630
rect 1177 31562 1297 31596
rect 1177 31528 1221 31562
rect 1255 31528 1297 31562
rect 1177 31494 1297 31528
rect 1177 31460 1221 31494
rect 1255 31460 1297 31494
rect 1177 31426 1297 31460
rect 1177 31392 1221 31426
rect 1255 31392 1297 31426
rect 1177 31358 1297 31392
rect 1177 31324 1221 31358
rect 1255 31324 1297 31358
rect 1177 31290 1297 31324
rect 1177 31256 1221 31290
rect 1255 31256 1297 31290
rect 1177 31222 1297 31256
rect 1177 31188 1221 31222
rect 1255 31188 1297 31222
rect 1177 31154 1297 31188
rect 1177 31120 1221 31154
rect 1255 31120 1297 31154
rect 1177 31086 1297 31120
rect 1177 31052 1221 31086
rect 1255 31052 1297 31086
rect 1177 31018 1297 31052
rect 1177 30984 1221 31018
rect 1255 30984 1297 31018
rect 1177 30950 1297 30984
rect 1177 30916 1221 30950
rect 1255 30916 1297 30950
rect 1177 30882 1297 30916
rect 1177 30848 1221 30882
rect 1255 30848 1297 30882
rect 1177 30814 1297 30848
rect 1177 30780 1221 30814
rect 1255 30780 1297 30814
rect 1177 30746 1297 30780
rect 1177 30712 1221 30746
rect 1255 30712 1297 30746
rect 1177 30678 1297 30712
rect 1177 30644 1221 30678
rect 1255 30644 1297 30678
rect 1177 30610 1297 30644
rect 1177 30576 1221 30610
rect 1255 30576 1297 30610
rect 1177 30542 1297 30576
rect 1177 30508 1221 30542
rect 1255 30508 1297 30542
rect 1177 30474 1297 30508
rect 1177 30440 1221 30474
rect 1255 30440 1297 30474
rect 1177 30406 1297 30440
rect 1177 30372 1221 30406
rect 1255 30372 1297 30406
rect 1177 30338 1297 30372
rect 1177 30304 1221 30338
rect 1255 30304 1297 30338
rect 1177 30270 1297 30304
rect 1177 30236 1221 30270
rect 1255 30236 1297 30270
rect 1177 30202 1297 30236
rect 1177 30168 1221 30202
rect 1255 30168 1297 30202
rect 1177 30134 1297 30168
rect 1177 30100 1221 30134
rect 1255 30100 1297 30134
rect 1177 30066 1297 30100
rect 1177 30032 1221 30066
rect 1255 30032 1297 30066
rect 1177 29998 1297 30032
rect 1177 29964 1221 29998
rect 1255 29964 1297 29998
rect 1177 29930 1297 29964
rect 1177 29896 1221 29930
rect 1255 29896 1297 29930
rect 1177 29862 1297 29896
rect 1177 29828 1221 29862
rect 1255 29828 1297 29862
rect 1177 29794 1297 29828
rect 1177 29760 1221 29794
rect 1255 29760 1297 29794
rect 1177 29726 1297 29760
rect 1177 29692 1221 29726
rect 1255 29692 1297 29726
rect 1177 29658 1297 29692
rect 1177 29624 1221 29658
rect 1255 29624 1297 29658
rect 1177 29590 1297 29624
rect 1177 29556 1221 29590
rect 1255 29556 1297 29590
rect 1177 29522 1297 29556
rect 1177 29488 1221 29522
rect 1255 29488 1297 29522
rect 1177 29454 1297 29488
rect 1177 29420 1221 29454
rect 1255 29420 1297 29454
rect 1177 29386 1297 29420
rect 1177 29352 1221 29386
rect 1255 29352 1297 29386
rect 1177 29318 1297 29352
rect 1177 29284 1221 29318
rect 1255 29284 1297 29318
rect 1177 29250 1297 29284
rect 1177 29216 1221 29250
rect 1255 29216 1297 29250
rect 1177 29182 1297 29216
rect 1177 29148 1221 29182
rect 1255 29148 1297 29182
rect 1177 29114 1297 29148
rect 1177 29080 1221 29114
rect 1255 29080 1297 29114
rect 1177 29046 1297 29080
rect 1177 29012 1221 29046
rect 1255 29012 1297 29046
rect 1177 28978 1297 29012
rect 1177 28944 1221 28978
rect 1255 28944 1297 28978
rect 1177 28910 1297 28944
rect 1177 28876 1221 28910
rect 1255 28876 1297 28910
rect 1177 28842 1297 28876
rect 1177 28808 1221 28842
rect 1255 28808 1297 28842
rect 1177 28774 1297 28808
rect 1177 28740 1221 28774
rect 1255 28740 1297 28774
rect 1177 28706 1297 28740
rect 1177 28672 1221 28706
rect 1255 28672 1297 28706
rect 1177 28638 1297 28672
rect 1177 28604 1221 28638
rect 1255 28604 1297 28638
rect 1177 28570 1297 28604
rect 1177 28536 1221 28570
rect 1255 28536 1297 28570
rect 1177 28502 1297 28536
rect 1177 28468 1221 28502
rect 1255 28468 1297 28502
rect 1177 28434 1297 28468
rect 1177 28400 1221 28434
rect 1255 28400 1297 28434
rect 1177 28366 1297 28400
rect 1177 28332 1221 28366
rect 1255 28332 1297 28366
rect 1177 28298 1297 28332
rect 1177 28264 1221 28298
rect 1255 28264 1297 28298
rect 1177 28230 1297 28264
rect 1177 28196 1221 28230
rect 1255 28196 1297 28230
rect 1177 28162 1297 28196
rect 1177 28128 1221 28162
rect 1255 28128 1297 28162
rect 1177 28094 1297 28128
rect 1177 28060 1221 28094
rect 1255 28060 1297 28094
rect 1177 28026 1297 28060
rect 1177 27992 1221 28026
rect 1255 27992 1297 28026
rect 1177 27958 1297 27992
rect 1177 27924 1221 27958
rect 1255 27924 1297 27958
rect 1177 27890 1297 27924
rect 1177 27856 1221 27890
rect 1255 27856 1297 27890
rect 1177 27822 1297 27856
rect 1177 27788 1221 27822
rect 1255 27788 1297 27822
rect 1177 27754 1297 27788
rect 1177 27720 1221 27754
rect 1255 27720 1297 27754
rect 1177 27686 1297 27720
rect 1177 27652 1221 27686
rect 1255 27652 1297 27686
rect 1177 27618 1297 27652
rect 1177 27584 1221 27618
rect 1255 27584 1297 27618
rect 1177 27550 1297 27584
rect 1177 27516 1221 27550
rect 1255 27516 1297 27550
rect 1177 27482 1297 27516
rect 1177 27448 1221 27482
rect 1255 27448 1297 27482
rect 1177 27414 1297 27448
rect 1177 27380 1221 27414
rect 1255 27380 1297 27414
rect 1177 27346 1297 27380
rect 1177 27312 1221 27346
rect 1255 27312 1297 27346
rect 1177 27278 1297 27312
rect 1177 27244 1221 27278
rect 1255 27244 1297 27278
rect 1177 27210 1297 27244
rect 1177 27176 1221 27210
rect 1255 27176 1297 27210
rect 1177 27142 1297 27176
rect 1177 27108 1221 27142
rect 1255 27108 1297 27142
rect 1177 27074 1297 27108
rect 1177 27040 1221 27074
rect 1255 27040 1297 27074
rect 1177 27006 1297 27040
rect 1177 26972 1221 27006
rect 1255 26972 1297 27006
rect 1177 26938 1297 26972
rect 1177 26904 1221 26938
rect 1255 26904 1297 26938
rect 1177 26870 1297 26904
rect 1177 26836 1221 26870
rect 1255 26836 1297 26870
rect 1177 26802 1297 26836
rect 1177 26768 1221 26802
rect 1255 26768 1297 26802
rect 1177 26734 1297 26768
rect 1177 26700 1221 26734
rect 1255 26700 1297 26734
rect 1177 26666 1297 26700
rect 1177 26632 1221 26666
rect 1255 26632 1297 26666
rect 1177 26598 1297 26632
rect 1177 26564 1221 26598
rect 1255 26564 1297 26598
rect 1177 26530 1297 26564
rect 1177 26496 1221 26530
rect 1255 26496 1297 26530
rect 1177 26462 1297 26496
rect 1177 26428 1221 26462
rect 1255 26428 1297 26462
rect 1177 26394 1297 26428
rect 1177 26360 1221 26394
rect 1255 26360 1297 26394
rect 1177 26326 1297 26360
rect 1177 26292 1221 26326
rect 1255 26292 1297 26326
rect 1177 26258 1297 26292
rect 1177 26224 1221 26258
rect 1255 26224 1297 26258
rect 1177 26190 1297 26224
rect 1177 26156 1221 26190
rect 1255 26156 1297 26190
rect 1177 26122 1297 26156
rect 1177 26088 1221 26122
rect 1255 26088 1297 26122
rect 1177 26054 1297 26088
rect 1177 26020 1221 26054
rect 1255 26020 1297 26054
rect 1177 25986 1297 26020
rect 1177 25952 1221 25986
rect 1255 25952 1297 25986
rect 1177 25918 1297 25952
rect 1177 25884 1221 25918
rect 1255 25884 1297 25918
rect 1177 25850 1297 25884
rect 1177 25816 1221 25850
rect 1255 25816 1297 25850
rect 1177 25782 1297 25816
rect 1177 25748 1221 25782
rect 1255 25748 1297 25782
rect 1177 25714 1297 25748
rect 1177 25680 1221 25714
rect 1255 25680 1297 25714
rect 1177 25646 1297 25680
rect 1177 25612 1221 25646
rect 1255 25612 1297 25646
rect 1177 25578 1297 25612
rect 1177 25544 1221 25578
rect 1255 25544 1297 25578
rect 1177 25510 1297 25544
rect 1177 25476 1221 25510
rect 1255 25476 1297 25510
rect 1177 25442 1297 25476
rect 1177 25408 1221 25442
rect 1255 25408 1297 25442
rect 1177 25374 1297 25408
rect 1177 25340 1221 25374
rect 1255 25340 1297 25374
rect 1177 25306 1297 25340
rect 1177 25272 1221 25306
rect 1255 25272 1297 25306
rect 1177 25238 1297 25272
rect 1177 25204 1221 25238
rect 1255 25204 1297 25238
rect 1177 25170 1297 25204
rect 1177 25136 1221 25170
rect 1255 25136 1297 25170
rect 1177 25102 1297 25136
rect 1177 25068 1221 25102
rect 1255 25068 1297 25102
rect 1177 25034 1297 25068
rect 1177 25000 1221 25034
rect 1255 25000 1297 25034
rect 1177 24966 1297 25000
rect 1177 24932 1221 24966
rect 1255 24932 1297 24966
rect 1177 24898 1297 24932
rect 1177 24864 1221 24898
rect 1255 24864 1297 24898
rect 1177 24830 1297 24864
rect 1177 24796 1221 24830
rect 1255 24796 1297 24830
rect 1177 24762 1297 24796
rect 1177 24728 1221 24762
rect 1255 24728 1297 24762
rect 1177 24694 1297 24728
rect 1177 24660 1221 24694
rect 1255 24660 1297 24694
rect 1177 24626 1297 24660
rect 1177 24592 1221 24626
rect 1255 24592 1297 24626
rect 1177 24558 1297 24592
rect 1177 24524 1221 24558
rect 1255 24524 1297 24558
rect 1177 24490 1297 24524
rect 1177 24456 1221 24490
rect 1255 24456 1297 24490
rect 1177 24422 1297 24456
rect 1177 24388 1221 24422
rect 1255 24388 1297 24422
rect 1177 24354 1297 24388
rect 1177 24320 1221 24354
rect 1255 24320 1297 24354
rect 1177 24286 1297 24320
rect 1177 24252 1221 24286
rect 1255 24252 1297 24286
rect 1177 24218 1297 24252
rect 1177 24184 1221 24218
rect 1255 24184 1297 24218
rect 1177 24150 1297 24184
rect 1177 24116 1221 24150
rect 1255 24116 1297 24150
rect 1177 24082 1297 24116
rect 1177 24048 1221 24082
rect 1255 24048 1297 24082
rect 1177 24014 1297 24048
rect 1177 23980 1221 24014
rect 1255 23980 1297 24014
rect 1177 23946 1297 23980
rect 1177 23912 1221 23946
rect 1255 23912 1297 23946
rect 1177 23878 1297 23912
rect 1177 23844 1221 23878
rect 1255 23844 1297 23878
rect 1177 23810 1297 23844
rect 1177 23776 1221 23810
rect 1255 23776 1297 23810
rect 1177 23742 1297 23776
rect 1177 23708 1221 23742
rect 1255 23708 1297 23742
rect 1177 23674 1297 23708
rect 1177 23640 1221 23674
rect 1255 23640 1297 23674
rect 1177 23606 1297 23640
rect 1177 23572 1221 23606
rect 1255 23572 1297 23606
rect 1177 23538 1297 23572
rect 1177 23504 1221 23538
rect 1255 23504 1297 23538
rect 1177 23470 1297 23504
rect 1177 23436 1221 23470
rect 1255 23436 1297 23470
rect 1177 23402 1297 23436
rect 1177 23368 1221 23402
rect 1255 23368 1297 23402
rect 1177 23334 1297 23368
rect 1177 23300 1221 23334
rect 1255 23300 1297 23334
rect 1177 23266 1297 23300
rect 1177 23232 1221 23266
rect 1255 23232 1297 23266
rect 1177 23198 1297 23232
rect 1177 23164 1221 23198
rect 1255 23164 1297 23198
rect 1177 23130 1297 23164
rect 1177 23096 1221 23130
rect 1255 23096 1297 23130
rect 1177 23062 1297 23096
rect 1177 23028 1221 23062
rect 1255 23028 1297 23062
rect 1177 22994 1297 23028
rect 1177 22960 1221 22994
rect 1255 22960 1297 22994
rect 1177 22926 1297 22960
rect 1177 22892 1221 22926
rect 1255 22892 1297 22926
rect 1177 22858 1297 22892
rect 1177 22824 1221 22858
rect 1255 22824 1297 22858
rect 1177 22790 1297 22824
rect 1177 22756 1221 22790
rect 1255 22756 1297 22790
rect 1177 22722 1297 22756
rect 1177 22688 1221 22722
rect 1255 22688 1297 22722
rect 1177 22654 1297 22688
rect 1177 22620 1221 22654
rect 1255 22620 1297 22654
rect 1177 22586 1297 22620
rect 1177 22552 1221 22586
rect 1255 22552 1297 22586
rect 1177 22518 1297 22552
rect 1177 22484 1221 22518
rect 1255 22484 1297 22518
rect 1177 22450 1297 22484
rect 1177 22416 1221 22450
rect 1255 22416 1297 22450
rect 1177 22382 1297 22416
rect 1177 22348 1221 22382
rect 1255 22348 1297 22382
rect 1177 22314 1297 22348
rect 1177 22280 1221 22314
rect 1255 22280 1297 22314
rect 1177 22246 1297 22280
rect 1177 22212 1221 22246
rect 1255 22212 1297 22246
rect 1177 22178 1297 22212
rect 1177 22144 1221 22178
rect 1255 22144 1297 22178
rect 1177 22110 1297 22144
rect 1177 22076 1221 22110
rect 1255 22076 1297 22110
rect 1177 22042 1297 22076
rect 1177 22008 1221 22042
rect 1255 22008 1297 22042
rect 1177 21974 1297 22008
rect 1177 21940 1221 21974
rect 1255 21940 1297 21974
rect 1177 21906 1297 21940
rect 1177 21872 1221 21906
rect 1255 21872 1297 21906
rect 1177 21838 1297 21872
rect 1177 21804 1221 21838
rect 1255 21804 1297 21838
rect 1177 21770 1297 21804
rect 1177 21736 1221 21770
rect 1255 21736 1297 21770
rect 1177 21702 1297 21736
rect 1177 21668 1221 21702
rect 1255 21668 1297 21702
rect 1177 21634 1297 21668
rect 1177 21600 1221 21634
rect 1255 21600 1297 21634
rect 1177 21566 1297 21600
rect 1177 21532 1221 21566
rect 1255 21532 1297 21566
rect 1177 21498 1297 21532
rect 1177 21464 1221 21498
rect 1255 21464 1297 21498
rect 1177 21430 1297 21464
rect 1177 21396 1221 21430
rect 1255 21396 1297 21430
rect 1177 21362 1297 21396
rect 1177 21328 1221 21362
rect 1255 21328 1297 21362
rect 1177 21294 1297 21328
rect 1177 21260 1221 21294
rect 1255 21260 1297 21294
rect 1177 21226 1297 21260
rect 1177 21192 1221 21226
rect 1255 21192 1297 21226
rect 1177 21158 1297 21192
rect 1177 21124 1221 21158
rect 1255 21124 1297 21158
rect 1177 21090 1297 21124
rect 1177 21056 1221 21090
rect 1255 21056 1297 21090
rect 1177 21022 1297 21056
rect 1177 20988 1221 21022
rect 1255 20988 1297 21022
rect 1177 20954 1297 20988
rect 1177 20920 1221 20954
rect 1255 20920 1297 20954
rect 1177 20886 1297 20920
rect 1177 20852 1221 20886
rect 1255 20852 1297 20886
rect 1177 20818 1297 20852
rect 1177 20784 1221 20818
rect 1255 20784 1297 20818
rect 1177 20750 1297 20784
rect 1177 20716 1221 20750
rect 1255 20716 1297 20750
rect 1177 20682 1297 20716
rect 1177 20648 1221 20682
rect 1255 20648 1297 20682
rect 1177 20614 1297 20648
rect 1177 20580 1221 20614
rect 1255 20580 1297 20614
rect 1177 20546 1297 20580
rect 1177 20512 1221 20546
rect 1255 20512 1297 20546
rect 1177 20478 1297 20512
rect 1177 20444 1221 20478
rect 1255 20444 1297 20478
rect 1177 20410 1297 20444
rect 1177 20376 1221 20410
rect 1255 20376 1297 20410
rect 1177 20342 1297 20376
rect 1177 20308 1221 20342
rect 1255 20308 1297 20342
rect 1177 20274 1297 20308
rect 1177 20240 1221 20274
rect 1255 20240 1297 20274
rect 1177 20206 1297 20240
rect 1177 20172 1221 20206
rect 1255 20172 1297 20206
rect 1177 20138 1297 20172
rect 1177 20104 1221 20138
rect 1255 20104 1297 20138
rect 1177 20070 1297 20104
rect 1177 20036 1221 20070
rect 1255 20036 1297 20070
rect 1177 20002 1297 20036
rect 1177 19968 1221 20002
rect 1255 19968 1297 20002
rect 1177 19934 1297 19968
rect 1177 19900 1221 19934
rect 1255 19900 1297 19934
rect 1177 19866 1297 19900
rect 1177 19832 1221 19866
rect 1255 19832 1297 19866
rect 1177 19798 1297 19832
rect 1177 19764 1221 19798
rect 1255 19764 1297 19798
rect 1177 19730 1297 19764
rect 1177 19696 1221 19730
rect 1255 19696 1297 19730
rect 1177 19662 1297 19696
rect 1177 19628 1221 19662
rect 1255 19628 1297 19662
rect 1177 19594 1297 19628
rect 1177 19560 1221 19594
rect 1255 19560 1297 19594
rect 1177 19526 1297 19560
rect 1177 19492 1221 19526
rect 1255 19492 1297 19526
rect 1177 19458 1297 19492
rect 1177 19424 1221 19458
rect 1255 19424 1297 19458
rect 1177 19390 1297 19424
rect 1177 19356 1221 19390
rect 1255 19356 1297 19390
rect 1177 19322 1297 19356
rect 1177 19288 1221 19322
rect 1255 19288 1297 19322
rect 1177 19254 1297 19288
rect 1177 19220 1221 19254
rect 1255 19220 1297 19254
rect 1177 19186 1297 19220
rect 1177 19152 1221 19186
rect 1255 19152 1297 19186
rect 1177 19118 1297 19152
rect 1177 19084 1221 19118
rect 1255 19084 1297 19118
rect 1177 19050 1297 19084
rect 1177 19016 1221 19050
rect 1255 19016 1297 19050
rect 1177 18982 1297 19016
rect 1177 18948 1221 18982
rect 1255 18948 1297 18982
rect 1177 18914 1297 18948
rect 1177 18880 1221 18914
rect 1255 18880 1297 18914
rect 1177 18846 1297 18880
rect 1177 18812 1221 18846
rect 1255 18812 1297 18846
rect 1177 18778 1297 18812
rect 1177 18744 1221 18778
rect 1255 18744 1297 18778
rect 1177 18710 1297 18744
rect 1177 18676 1221 18710
rect 1255 18676 1297 18710
rect 1177 18642 1297 18676
rect 1177 18608 1221 18642
rect 1255 18608 1297 18642
rect 1177 18574 1297 18608
rect 1177 18540 1221 18574
rect 1255 18540 1297 18574
rect 1177 18506 1297 18540
rect 1177 18472 1221 18506
rect 1255 18472 1297 18506
rect 1177 18438 1297 18472
rect 1177 18404 1221 18438
rect 1255 18404 1297 18438
rect 1177 18370 1297 18404
rect 1177 18336 1221 18370
rect 1255 18336 1297 18370
rect 1177 18302 1297 18336
rect 1177 18268 1221 18302
rect 1255 18268 1297 18302
rect 1177 18234 1297 18268
rect 1177 18200 1221 18234
rect 1255 18200 1297 18234
rect 1177 18166 1297 18200
rect 1177 18132 1221 18166
rect 1255 18132 1297 18166
rect 1177 18098 1297 18132
rect 1177 18064 1221 18098
rect 1255 18064 1297 18098
rect 1177 18030 1297 18064
rect 1177 17996 1221 18030
rect 1255 17996 1297 18030
rect 1177 17962 1297 17996
rect 1177 17928 1221 17962
rect 1255 17928 1297 17962
rect 1177 17894 1297 17928
rect 1177 17860 1221 17894
rect 1255 17860 1297 17894
rect 1177 17826 1297 17860
rect 1177 17792 1221 17826
rect 1255 17792 1297 17826
rect 1177 17758 1297 17792
rect 1177 17724 1221 17758
rect 1255 17724 1297 17758
rect 1177 17690 1297 17724
rect 1177 17656 1221 17690
rect 1255 17656 1297 17690
rect 1177 17622 1297 17656
rect 1177 17588 1221 17622
rect 1255 17588 1297 17622
rect 1177 17554 1297 17588
rect 1177 17520 1221 17554
rect 1255 17520 1297 17554
rect 1177 17486 1297 17520
rect 1177 17452 1221 17486
rect 1255 17452 1297 17486
rect 1177 17418 1297 17452
rect 1177 17384 1221 17418
rect 1255 17384 1297 17418
rect 1177 17350 1297 17384
rect 1177 17316 1221 17350
rect 1255 17316 1297 17350
rect 1177 17282 1297 17316
rect 1177 17248 1221 17282
rect 1255 17248 1297 17282
rect 1177 17214 1297 17248
rect 1177 17180 1221 17214
rect 1255 17180 1297 17214
rect 1177 17146 1297 17180
rect 1177 17112 1221 17146
rect 1255 17112 1297 17146
rect 1177 17078 1297 17112
rect 1177 17044 1221 17078
rect 1255 17044 1297 17078
rect 1177 17010 1297 17044
rect 1177 16976 1221 17010
rect 1255 16976 1297 17010
rect 1177 16942 1297 16976
rect 1177 16908 1221 16942
rect 1255 16908 1297 16942
rect 1177 16874 1297 16908
rect 1177 16840 1221 16874
rect 1255 16840 1297 16874
rect 1177 16806 1297 16840
rect 1177 16772 1221 16806
rect 1255 16772 1297 16806
rect 1177 16738 1297 16772
rect 1177 16704 1221 16738
rect 1255 16704 1297 16738
rect 1177 16670 1297 16704
rect 1177 16636 1221 16670
rect 1255 16636 1297 16670
rect 1177 16602 1297 16636
rect 1177 16568 1221 16602
rect 1255 16568 1297 16602
rect 1177 16534 1297 16568
rect 1177 16500 1221 16534
rect 1255 16500 1297 16534
rect 1177 16466 1297 16500
rect 1177 16432 1221 16466
rect 1255 16432 1297 16466
rect 1177 16398 1297 16432
rect 1177 16364 1221 16398
rect 1255 16364 1297 16398
rect 1177 16330 1297 16364
rect 1177 16296 1221 16330
rect 1255 16296 1297 16330
rect 1177 16262 1297 16296
rect 1177 16228 1221 16262
rect 1255 16228 1297 16262
rect 1177 16194 1297 16228
rect 1177 16160 1221 16194
rect 1255 16160 1297 16194
rect 1177 16126 1297 16160
rect 1177 16092 1221 16126
rect 1255 16092 1297 16126
rect 1177 16058 1297 16092
rect 1177 16024 1221 16058
rect 1255 16024 1297 16058
rect 1177 15990 1297 16024
rect 1177 15956 1221 15990
rect 1255 15956 1297 15990
rect 1177 15922 1297 15956
rect 1177 15888 1221 15922
rect 1255 15888 1297 15922
rect 1177 15854 1297 15888
rect 1177 15820 1221 15854
rect 1255 15820 1297 15854
rect 1177 15786 1297 15820
rect 1177 15752 1221 15786
rect 1255 15752 1297 15786
rect 1177 15718 1297 15752
rect 1177 15684 1221 15718
rect 1255 15684 1297 15718
rect 1177 15650 1297 15684
rect 1177 15616 1221 15650
rect 1255 15616 1297 15650
rect 1177 15582 1297 15616
rect 1177 15548 1221 15582
rect 1255 15548 1297 15582
rect 1177 15514 1297 15548
rect 1177 15480 1221 15514
rect 1255 15480 1297 15514
rect 1177 15446 1297 15480
rect 1177 15412 1221 15446
rect 1255 15412 1297 15446
rect 1177 15378 1297 15412
rect 1177 15344 1221 15378
rect 1255 15344 1297 15378
rect 1177 15310 1297 15344
rect 1177 15276 1221 15310
rect 1255 15276 1297 15310
rect 1177 15242 1297 15276
rect 1177 15208 1221 15242
rect 1255 15208 1297 15242
rect 1177 15174 1297 15208
rect 1177 15140 1221 15174
rect 1255 15140 1297 15174
rect 1177 15106 1297 15140
rect 1177 15072 1221 15106
rect 1255 15072 1297 15106
rect 1177 15038 1297 15072
rect 1177 15004 1221 15038
rect 1255 15004 1297 15038
rect 1177 14970 1297 15004
rect 1177 14936 1221 14970
rect 1255 14936 1297 14970
rect 1177 14902 1297 14936
rect 1177 14868 1221 14902
rect 1255 14868 1297 14902
rect 1177 14834 1297 14868
rect 1177 14800 1221 14834
rect 1255 14800 1297 14834
rect 1177 14766 1297 14800
rect 1177 14732 1221 14766
rect 1255 14732 1297 14766
rect 1177 14698 1297 14732
rect 1177 14664 1221 14698
rect 1255 14664 1297 14698
rect 1177 14630 1297 14664
rect 1177 14596 1221 14630
rect 1255 14596 1297 14630
rect 1177 14562 1297 14596
rect 1177 14528 1221 14562
rect 1255 14528 1297 14562
rect 1177 14494 1297 14528
rect 1177 14460 1221 14494
rect 1255 14460 1297 14494
rect 1177 14426 1297 14460
rect 1177 14392 1221 14426
rect 1255 14392 1297 14426
rect 1177 14358 1297 14392
rect 1177 14324 1221 14358
rect 1255 14324 1297 14358
rect 1177 14290 1297 14324
rect 1177 14256 1221 14290
rect 1255 14256 1297 14290
rect 1177 14222 1297 14256
rect 1177 14188 1221 14222
rect 1255 14188 1297 14222
rect 1177 14154 1297 14188
rect 1177 14120 1221 14154
rect 1255 14120 1297 14154
rect 1177 14086 1297 14120
rect 1177 14052 1221 14086
rect 1255 14052 1297 14086
rect 1177 14018 1297 14052
rect 1177 13984 1221 14018
rect 1255 13984 1297 14018
rect 1177 13950 1297 13984
rect 1177 13916 1221 13950
rect 1255 13916 1297 13950
rect 1177 13882 1297 13916
rect 1177 13848 1221 13882
rect 1255 13848 1297 13882
rect 1177 13814 1297 13848
rect 1177 13780 1221 13814
rect 1255 13780 1297 13814
rect 1177 13746 1297 13780
rect 1177 13712 1221 13746
rect 1255 13712 1297 13746
rect 1177 13678 1297 13712
rect 1177 13644 1221 13678
rect 1255 13644 1297 13678
rect 1177 13610 1297 13644
rect 1177 13576 1221 13610
rect 1255 13576 1297 13610
rect 1177 13542 1297 13576
rect 1177 13508 1221 13542
rect 1255 13508 1297 13542
rect 1177 13474 1297 13508
rect 1177 13440 1221 13474
rect 1255 13440 1297 13474
rect 1177 13406 1297 13440
rect 1177 13372 1221 13406
rect 1255 13372 1297 13406
rect 1177 13338 1297 13372
rect 1177 13304 1221 13338
rect 1255 13304 1297 13338
rect 1177 13270 1297 13304
rect 1177 13236 1221 13270
rect 1255 13236 1297 13270
rect 1177 13202 1297 13236
rect 1177 13168 1221 13202
rect 1255 13168 1297 13202
rect 1177 13134 1297 13168
rect 1177 13100 1221 13134
rect 1255 13100 1297 13134
rect 1177 13066 1297 13100
rect 1177 13032 1221 13066
rect 1255 13032 1297 13066
rect 1177 12998 1297 13032
rect 1177 12964 1221 12998
rect 1255 12964 1297 12998
rect 1177 12930 1297 12964
rect 1177 12896 1221 12930
rect 1255 12896 1297 12930
rect 1177 12862 1297 12896
rect 1177 12828 1221 12862
rect 1255 12828 1297 12862
rect 1177 12794 1297 12828
rect 1177 12760 1221 12794
rect 1255 12760 1297 12794
rect 1177 12726 1297 12760
rect 1177 12692 1221 12726
rect 1255 12692 1297 12726
rect 1177 12658 1297 12692
rect 1177 12624 1221 12658
rect 1255 12624 1297 12658
rect 1177 12590 1297 12624
rect 1177 12556 1221 12590
rect 1255 12556 1297 12590
rect 1177 12522 1297 12556
rect 1177 12488 1221 12522
rect 1255 12488 1297 12522
rect 1177 12454 1297 12488
rect 1177 12420 1221 12454
rect 1255 12420 1297 12454
rect 1177 12386 1297 12420
rect 1177 12352 1221 12386
rect 1255 12352 1297 12386
rect 1177 12318 1297 12352
rect 1177 12284 1221 12318
rect 1255 12284 1297 12318
rect 1177 12250 1297 12284
rect 1177 12216 1221 12250
rect 1255 12216 1297 12250
rect 1177 12182 1297 12216
rect 1177 12148 1221 12182
rect 1255 12148 1297 12182
rect 1177 12114 1297 12148
rect 1177 12080 1221 12114
rect 1255 12080 1297 12114
rect 1177 12046 1297 12080
rect 1177 12012 1221 12046
rect 1255 12012 1297 12046
rect 1177 11978 1297 12012
rect 1177 11944 1221 11978
rect 1255 11944 1297 11978
rect 1177 11910 1297 11944
rect 1177 11876 1221 11910
rect 1255 11876 1297 11910
rect 1177 11842 1297 11876
rect 1177 11808 1221 11842
rect 1255 11808 1297 11842
rect 1177 11774 1297 11808
rect 1177 11740 1221 11774
rect 1255 11740 1297 11774
rect 1177 11706 1297 11740
rect 1177 11672 1221 11706
rect 1255 11672 1297 11706
rect 1177 11638 1297 11672
rect 1177 11604 1221 11638
rect 1255 11604 1297 11638
rect 1177 11570 1297 11604
rect 1177 11536 1221 11570
rect 1255 11536 1297 11570
rect 1177 11502 1297 11536
rect 1177 11468 1221 11502
rect 1255 11468 1297 11502
rect 1177 11434 1297 11468
rect 1177 11400 1221 11434
rect 1255 11400 1297 11434
rect 1177 11366 1297 11400
rect 1177 11332 1221 11366
rect 1255 11332 1297 11366
rect 1177 11298 1297 11332
rect 1177 11264 1221 11298
rect 1255 11264 1297 11298
rect 1177 11230 1297 11264
rect 1177 11196 1221 11230
rect 1255 11196 1297 11230
rect 1177 11162 1297 11196
rect 1177 11128 1221 11162
rect 1255 11128 1297 11162
rect 1177 11094 1297 11128
rect 1177 11060 1221 11094
rect 1255 11060 1297 11094
rect 1177 11026 1297 11060
rect 1177 10992 1221 11026
rect 1255 10992 1297 11026
rect 1177 10958 1297 10992
rect 1177 10924 1221 10958
rect 1255 10924 1297 10958
rect 1177 10890 1297 10924
rect 1177 10856 1221 10890
rect 1255 10856 1297 10890
rect 1177 10822 1297 10856
rect 1177 10788 1221 10822
rect 1255 10788 1297 10822
rect 1177 10754 1297 10788
rect 1177 10720 1221 10754
rect 1255 10720 1297 10754
rect 1177 10686 1297 10720
rect 1177 10652 1221 10686
rect 1255 10652 1297 10686
rect 1177 10618 1297 10652
rect 1177 10584 1221 10618
rect 1255 10584 1297 10618
rect 1177 10550 1297 10584
rect 1177 10516 1221 10550
rect 1255 10516 1297 10550
rect 1177 10482 1297 10516
rect 1177 10448 1221 10482
rect 1255 10448 1297 10482
rect 1177 10414 1297 10448
rect 1177 10380 1221 10414
rect 1255 10380 1297 10414
rect 1177 10334 1297 10380
rect 13697 34490 13817 34564
rect 13697 34456 13739 34490
rect 13773 34456 13817 34490
rect 13697 34422 13817 34456
rect 13697 34388 13739 34422
rect 13773 34388 13817 34422
rect 13697 34354 13817 34388
rect 13697 34320 13739 34354
rect 13773 34320 13817 34354
rect 13697 34286 13817 34320
rect 13697 34252 13739 34286
rect 13773 34252 13817 34286
rect 13697 34218 13817 34252
rect 13697 34184 13739 34218
rect 13773 34184 13817 34218
rect 13697 34150 13817 34184
rect 13697 34116 13739 34150
rect 13773 34116 13817 34150
rect 13697 34082 13817 34116
rect 13697 34048 13739 34082
rect 13773 34048 13817 34082
rect 13697 34014 13817 34048
rect 13697 33980 13739 34014
rect 13773 33980 13817 34014
rect 13697 33946 13817 33980
rect 13697 33912 13739 33946
rect 13773 33912 13817 33946
rect 13697 33878 13817 33912
rect 13697 33844 13739 33878
rect 13773 33844 13817 33878
rect 13697 33810 13817 33844
rect 13697 33776 13739 33810
rect 13773 33776 13817 33810
rect 13697 33742 13817 33776
rect 13697 33708 13739 33742
rect 13773 33708 13817 33742
rect 13697 33674 13817 33708
rect 13697 33640 13739 33674
rect 13773 33640 13817 33674
rect 13697 33606 13817 33640
rect 13697 33572 13739 33606
rect 13773 33572 13817 33606
rect 13697 33538 13817 33572
rect 13697 33504 13739 33538
rect 13773 33504 13817 33538
rect 13697 33470 13817 33504
rect 13697 33436 13739 33470
rect 13773 33436 13817 33470
rect 13697 33402 13817 33436
rect 13697 33368 13739 33402
rect 13773 33368 13817 33402
rect 13697 33334 13817 33368
rect 13697 33300 13739 33334
rect 13773 33300 13817 33334
rect 13697 33266 13817 33300
rect 13697 33232 13739 33266
rect 13773 33232 13817 33266
rect 13697 33198 13817 33232
rect 13697 33164 13739 33198
rect 13773 33164 13817 33198
rect 13697 33130 13817 33164
rect 13697 33096 13739 33130
rect 13773 33096 13817 33130
rect 13697 33062 13817 33096
rect 13697 33028 13739 33062
rect 13773 33028 13817 33062
rect 13697 32994 13817 33028
rect 13697 32960 13739 32994
rect 13773 32960 13817 32994
rect 13697 32926 13817 32960
rect 13697 32892 13739 32926
rect 13773 32892 13817 32926
rect 13697 32858 13817 32892
rect 13697 32824 13739 32858
rect 13773 32824 13817 32858
rect 13697 32790 13817 32824
rect 13697 32756 13739 32790
rect 13773 32756 13817 32790
rect 13697 32722 13817 32756
rect 13697 32688 13739 32722
rect 13773 32688 13817 32722
rect 13697 32654 13817 32688
rect 13697 32620 13739 32654
rect 13773 32620 13817 32654
rect 13697 32586 13817 32620
rect 13697 32552 13739 32586
rect 13773 32552 13817 32586
rect 13697 32518 13817 32552
rect 13697 32484 13739 32518
rect 13773 32484 13817 32518
rect 13697 32450 13817 32484
rect 13697 32416 13739 32450
rect 13773 32416 13817 32450
rect 13697 32382 13817 32416
rect 13697 32348 13739 32382
rect 13773 32348 13817 32382
rect 13697 32314 13817 32348
rect 13697 32280 13739 32314
rect 13773 32280 13817 32314
rect 13697 32246 13817 32280
rect 13697 32212 13739 32246
rect 13773 32212 13817 32246
rect 13697 32178 13817 32212
rect 13697 32144 13739 32178
rect 13773 32144 13817 32178
rect 13697 32110 13817 32144
rect 13697 32076 13739 32110
rect 13773 32076 13817 32110
rect 13697 32042 13817 32076
rect 13697 32008 13739 32042
rect 13773 32008 13817 32042
rect 13697 31974 13817 32008
rect 13697 31940 13739 31974
rect 13773 31940 13817 31974
rect 13697 31906 13817 31940
rect 13697 31872 13739 31906
rect 13773 31872 13817 31906
rect 13697 31838 13817 31872
rect 13697 31804 13739 31838
rect 13773 31804 13817 31838
rect 13697 31770 13817 31804
rect 13697 31736 13739 31770
rect 13773 31736 13817 31770
rect 13697 31702 13817 31736
rect 13697 31668 13739 31702
rect 13773 31668 13817 31702
rect 13697 31634 13817 31668
rect 13697 31600 13739 31634
rect 13773 31600 13817 31634
rect 13697 31566 13817 31600
rect 13697 31532 13739 31566
rect 13773 31532 13817 31566
rect 13697 31498 13817 31532
rect 13697 31464 13739 31498
rect 13773 31464 13817 31498
rect 13697 31430 13817 31464
rect 13697 31396 13739 31430
rect 13773 31396 13817 31430
rect 13697 31362 13817 31396
rect 13697 31328 13739 31362
rect 13773 31328 13817 31362
rect 13697 31294 13817 31328
rect 13697 31260 13739 31294
rect 13773 31260 13817 31294
rect 13697 31226 13817 31260
rect 13697 31192 13739 31226
rect 13773 31192 13817 31226
rect 13697 31158 13817 31192
rect 13697 31124 13739 31158
rect 13773 31124 13817 31158
rect 13697 31090 13817 31124
rect 13697 31056 13739 31090
rect 13773 31056 13817 31090
rect 13697 31022 13817 31056
rect 13697 30988 13739 31022
rect 13773 30988 13817 31022
rect 13697 30954 13817 30988
rect 13697 30920 13739 30954
rect 13773 30920 13817 30954
rect 13697 30886 13817 30920
rect 13697 30852 13739 30886
rect 13773 30852 13817 30886
rect 13697 30818 13817 30852
rect 13697 30784 13739 30818
rect 13773 30784 13817 30818
rect 13697 30750 13817 30784
rect 13697 30716 13739 30750
rect 13773 30716 13817 30750
rect 13697 30682 13817 30716
rect 13697 30648 13739 30682
rect 13773 30648 13817 30682
rect 13697 30614 13817 30648
rect 13697 30580 13739 30614
rect 13773 30580 13817 30614
rect 13697 30546 13817 30580
rect 13697 30512 13739 30546
rect 13773 30512 13817 30546
rect 13697 30478 13817 30512
rect 13697 30444 13739 30478
rect 13773 30444 13817 30478
rect 13697 30410 13817 30444
rect 13697 30376 13739 30410
rect 13773 30376 13817 30410
rect 13697 30342 13817 30376
rect 13697 30308 13739 30342
rect 13773 30308 13817 30342
rect 13697 30274 13817 30308
rect 13697 30240 13739 30274
rect 13773 30240 13817 30274
rect 13697 30206 13817 30240
rect 13697 30172 13739 30206
rect 13773 30172 13817 30206
rect 13697 30138 13817 30172
rect 13697 30104 13739 30138
rect 13773 30104 13817 30138
rect 13697 30070 13817 30104
rect 13697 30036 13739 30070
rect 13773 30036 13817 30070
rect 13697 30002 13817 30036
rect 13697 29968 13739 30002
rect 13773 29968 13817 30002
rect 13697 29934 13817 29968
rect 13697 29900 13739 29934
rect 13773 29900 13817 29934
rect 13697 29866 13817 29900
rect 13697 29832 13739 29866
rect 13773 29832 13817 29866
rect 13697 29798 13817 29832
rect 13697 29764 13739 29798
rect 13773 29764 13817 29798
rect 13697 29730 13817 29764
rect 13697 29696 13739 29730
rect 13773 29696 13817 29730
rect 13697 29662 13817 29696
rect 13697 29628 13739 29662
rect 13773 29628 13817 29662
rect 13697 29594 13817 29628
rect 13697 29560 13739 29594
rect 13773 29560 13817 29594
rect 13697 29526 13817 29560
rect 13697 29492 13739 29526
rect 13773 29492 13817 29526
rect 13697 29458 13817 29492
rect 13697 29424 13739 29458
rect 13773 29424 13817 29458
rect 13697 29390 13817 29424
rect 13697 29356 13739 29390
rect 13773 29356 13817 29390
rect 13697 29322 13817 29356
rect 13697 29288 13739 29322
rect 13773 29288 13817 29322
rect 13697 29254 13817 29288
rect 13697 29220 13739 29254
rect 13773 29220 13817 29254
rect 13697 29186 13817 29220
rect 13697 29152 13739 29186
rect 13773 29152 13817 29186
rect 13697 29118 13817 29152
rect 13697 29084 13739 29118
rect 13773 29084 13817 29118
rect 13697 29050 13817 29084
rect 13697 29016 13739 29050
rect 13773 29016 13817 29050
rect 13697 28982 13817 29016
rect 13697 28948 13739 28982
rect 13773 28948 13817 28982
rect 13697 28914 13817 28948
rect 13697 28880 13739 28914
rect 13773 28880 13817 28914
rect 13697 28846 13817 28880
rect 13697 28812 13739 28846
rect 13773 28812 13817 28846
rect 13697 28778 13817 28812
rect 13697 28744 13739 28778
rect 13773 28744 13817 28778
rect 13697 28710 13817 28744
rect 13697 28676 13739 28710
rect 13773 28676 13817 28710
rect 13697 28642 13817 28676
rect 13697 28608 13739 28642
rect 13773 28608 13817 28642
rect 13697 28574 13817 28608
rect 13697 28540 13739 28574
rect 13773 28540 13817 28574
rect 13697 28506 13817 28540
rect 13697 28472 13739 28506
rect 13773 28472 13817 28506
rect 13697 28438 13817 28472
rect 13697 28404 13739 28438
rect 13773 28404 13817 28438
rect 13697 28370 13817 28404
rect 13697 28336 13739 28370
rect 13773 28336 13817 28370
rect 13697 28302 13817 28336
rect 13697 28268 13739 28302
rect 13773 28268 13817 28302
rect 13697 28234 13817 28268
rect 13697 28200 13739 28234
rect 13773 28200 13817 28234
rect 13697 28166 13817 28200
rect 13697 28132 13739 28166
rect 13773 28132 13817 28166
rect 13697 28098 13817 28132
rect 13697 28064 13739 28098
rect 13773 28064 13817 28098
rect 13697 28030 13817 28064
rect 13697 27996 13739 28030
rect 13773 27996 13817 28030
rect 13697 27962 13817 27996
rect 13697 27928 13739 27962
rect 13773 27928 13817 27962
rect 13697 27894 13817 27928
rect 13697 27860 13739 27894
rect 13773 27860 13817 27894
rect 13697 27826 13817 27860
rect 13697 27792 13739 27826
rect 13773 27792 13817 27826
rect 13697 27758 13817 27792
rect 13697 27724 13739 27758
rect 13773 27724 13817 27758
rect 13697 27690 13817 27724
rect 13697 27656 13739 27690
rect 13773 27656 13817 27690
rect 13697 27622 13817 27656
rect 13697 27588 13739 27622
rect 13773 27588 13817 27622
rect 13697 27554 13817 27588
rect 13697 27520 13739 27554
rect 13773 27520 13817 27554
rect 13697 27486 13817 27520
rect 13697 27452 13739 27486
rect 13773 27452 13817 27486
rect 13697 27418 13817 27452
rect 13697 27384 13739 27418
rect 13773 27384 13817 27418
rect 13697 27350 13817 27384
rect 13697 27316 13739 27350
rect 13773 27316 13817 27350
rect 13697 27282 13817 27316
rect 13697 27248 13739 27282
rect 13773 27248 13817 27282
rect 13697 27214 13817 27248
rect 13697 27180 13739 27214
rect 13773 27180 13817 27214
rect 13697 27146 13817 27180
rect 13697 27112 13739 27146
rect 13773 27112 13817 27146
rect 13697 27078 13817 27112
rect 13697 27044 13739 27078
rect 13773 27044 13817 27078
rect 13697 27010 13817 27044
rect 13697 26976 13739 27010
rect 13773 26976 13817 27010
rect 13697 26942 13817 26976
rect 13697 26908 13739 26942
rect 13773 26908 13817 26942
rect 13697 26874 13817 26908
rect 13697 26840 13739 26874
rect 13773 26840 13817 26874
rect 13697 26806 13817 26840
rect 13697 26772 13739 26806
rect 13773 26772 13817 26806
rect 13697 26738 13817 26772
rect 13697 26704 13739 26738
rect 13773 26704 13817 26738
rect 13697 26670 13817 26704
rect 13697 26636 13739 26670
rect 13773 26636 13817 26670
rect 13697 26602 13817 26636
rect 13697 26568 13739 26602
rect 13773 26568 13817 26602
rect 13697 26534 13817 26568
rect 13697 26500 13739 26534
rect 13773 26500 13817 26534
rect 13697 26466 13817 26500
rect 13697 26432 13739 26466
rect 13773 26432 13817 26466
rect 13697 26398 13817 26432
rect 13697 26364 13739 26398
rect 13773 26364 13817 26398
rect 13697 26330 13817 26364
rect 13697 26296 13739 26330
rect 13773 26296 13817 26330
rect 13697 26262 13817 26296
rect 13697 26228 13739 26262
rect 13773 26228 13817 26262
rect 13697 26194 13817 26228
rect 13697 26160 13739 26194
rect 13773 26160 13817 26194
rect 13697 26126 13817 26160
rect 13697 26092 13739 26126
rect 13773 26092 13817 26126
rect 13697 26058 13817 26092
rect 13697 26024 13739 26058
rect 13773 26024 13817 26058
rect 13697 25990 13817 26024
rect 13697 25956 13739 25990
rect 13773 25956 13817 25990
rect 13697 25922 13817 25956
rect 13697 25888 13739 25922
rect 13773 25888 13817 25922
rect 13697 25854 13817 25888
rect 13697 25820 13739 25854
rect 13773 25820 13817 25854
rect 13697 25786 13817 25820
rect 13697 25752 13739 25786
rect 13773 25752 13817 25786
rect 13697 25718 13817 25752
rect 13697 25684 13739 25718
rect 13773 25684 13817 25718
rect 13697 25650 13817 25684
rect 13697 25616 13739 25650
rect 13773 25616 13817 25650
rect 13697 25582 13817 25616
rect 13697 25548 13739 25582
rect 13773 25548 13817 25582
rect 13697 25514 13817 25548
rect 13697 25480 13739 25514
rect 13773 25480 13817 25514
rect 13697 25446 13817 25480
rect 13697 25412 13739 25446
rect 13773 25412 13817 25446
rect 13697 25378 13817 25412
rect 13697 25344 13739 25378
rect 13773 25344 13817 25378
rect 13697 25310 13817 25344
rect 13697 25276 13739 25310
rect 13773 25276 13817 25310
rect 13697 25242 13817 25276
rect 13697 25208 13739 25242
rect 13773 25208 13817 25242
rect 13697 25174 13817 25208
rect 13697 25140 13739 25174
rect 13773 25140 13817 25174
rect 13697 25106 13817 25140
rect 13697 25072 13739 25106
rect 13773 25072 13817 25106
rect 13697 25038 13817 25072
rect 13697 25004 13739 25038
rect 13773 25004 13817 25038
rect 13697 24970 13817 25004
rect 13697 24936 13739 24970
rect 13773 24936 13817 24970
rect 13697 24902 13817 24936
rect 13697 24868 13739 24902
rect 13773 24868 13817 24902
rect 13697 24834 13817 24868
rect 13697 24800 13739 24834
rect 13773 24800 13817 24834
rect 13697 24766 13817 24800
rect 13697 24732 13739 24766
rect 13773 24732 13817 24766
rect 13697 24698 13817 24732
rect 13697 24664 13739 24698
rect 13773 24664 13817 24698
rect 13697 24630 13817 24664
rect 13697 24596 13739 24630
rect 13773 24596 13817 24630
rect 13697 24562 13817 24596
rect 13697 24528 13739 24562
rect 13773 24528 13817 24562
rect 13697 24494 13817 24528
rect 13697 24460 13739 24494
rect 13773 24460 13817 24494
rect 13697 24426 13817 24460
rect 13697 24392 13739 24426
rect 13773 24392 13817 24426
rect 13697 24358 13817 24392
rect 13697 24324 13739 24358
rect 13773 24324 13817 24358
rect 13697 24290 13817 24324
rect 13697 24256 13739 24290
rect 13773 24256 13817 24290
rect 13697 24222 13817 24256
rect 13697 24188 13739 24222
rect 13773 24188 13817 24222
rect 13697 24154 13817 24188
rect 13697 24120 13739 24154
rect 13773 24120 13817 24154
rect 13697 24086 13817 24120
rect 13697 24052 13739 24086
rect 13773 24052 13817 24086
rect 13697 24018 13817 24052
rect 13697 23984 13739 24018
rect 13773 23984 13817 24018
rect 13697 23950 13817 23984
rect 13697 23916 13739 23950
rect 13773 23916 13817 23950
rect 13697 23882 13817 23916
rect 13697 23848 13739 23882
rect 13773 23848 13817 23882
rect 13697 23814 13817 23848
rect 13697 23780 13739 23814
rect 13773 23780 13817 23814
rect 13697 23746 13817 23780
rect 13697 23712 13739 23746
rect 13773 23712 13817 23746
rect 13697 23678 13817 23712
rect 13697 23644 13739 23678
rect 13773 23644 13817 23678
rect 13697 23610 13817 23644
rect 13697 23576 13739 23610
rect 13773 23576 13817 23610
rect 13697 23542 13817 23576
rect 13697 23508 13739 23542
rect 13773 23508 13817 23542
rect 13697 23474 13817 23508
rect 13697 23440 13739 23474
rect 13773 23440 13817 23474
rect 13697 23406 13817 23440
rect 13697 23372 13739 23406
rect 13773 23372 13817 23406
rect 13697 23338 13817 23372
rect 13697 23304 13739 23338
rect 13773 23304 13817 23338
rect 13697 23270 13817 23304
rect 13697 23236 13739 23270
rect 13773 23236 13817 23270
rect 13697 23202 13817 23236
rect 13697 23168 13739 23202
rect 13773 23168 13817 23202
rect 13697 23134 13817 23168
rect 13697 23100 13739 23134
rect 13773 23100 13817 23134
rect 13697 23066 13817 23100
rect 13697 23032 13739 23066
rect 13773 23032 13817 23066
rect 13697 22998 13817 23032
rect 13697 22964 13739 22998
rect 13773 22964 13817 22998
rect 13697 22930 13817 22964
rect 13697 22896 13739 22930
rect 13773 22896 13817 22930
rect 13697 22862 13817 22896
rect 13697 22828 13739 22862
rect 13773 22828 13817 22862
rect 13697 22794 13817 22828
rect 13697 22760 13739 22794
rect 13773 22760 13817 22794
rect 13697 22726 13817 22760
rect 13697 22692 13739 22726
rect 13773 22692 13817 22726
rect 13697 22658 13817 22692
rect 13697 22624 13739 22658
rect 13773 22624 13817 22658
rect 13697 22590 13817 22624
rect 13697 22556 13739 22590
rect 13773 22556 13817 22590
rect 13697 22522 13817 22556
rect 13697 22488 13739 22522
rect 13773 22488 13817 22522
rect 13697 22454 13817 22488
rect 13697 22420 13739 22454
rect 13773 22420 13817 22454
rect 13697 22386 13817 22420
rect 13697 22352 13739 22386
rect 13773 22352 13817 22386
rect 13697 22318 13817 22352
rect 13697 22284 13739 22318
rect 13773 22284 13817 22318
rect 13697 22250 13817 22284
rect 13697 22216 13739 22250
rect 13773 22216 13817 22250
rect 13697 22182 13817 22216
rect 13697 22148 13739 22182
rect 13773 22148 13817 22182
rect 13697 22114 13817 22148
rect 13697 22080 13739 22114
rect 13773 22080 13817 22114
rect 13697 22046 13817 22080
rect 13697 22012 13739 22046
rect 13773 22012 13817 22046
rect 13697 21978 13817 22012
rect 13697 21944 13739 21978
rect 13773 21944 13817 21978
rect 13697 21910 13817 21944
rect 13697 21876 13739 21910
rect 13773 21876 13817 21910
rect 13697 21842 13817 21876
rect 13697 21808 13739 21842
rect 13773 21808 13817 21842
rect 13697 21774 13817 21808
rect 13697 21740 13739 21774
rect 13773 21740 13817 21774
rect 13697 21706 13817 21740
rect 13697 21672 13739 21706
rect 13773 21672 13817 21706
rect 13697 21638 13817 21672
rect 13697 21604 13739 21638
rect 13773 21604 13817 21638
rect 13697 21570 13817 21604
rect 13697 21536 13739 21570
rect 13773 21536 13817 21570
rect 13697 21502 13817 21536
rect 13697 21468 13739 21502
rect 13773 21468 13817 21502
rect 13697 21434 13817 21468
rect 13697 21400 13739 21434
rect 13773 21400 13817 21434
rect 13697 21366 13817 21400
rect 13697 21332 13739 21366
rect 13773 21332 13817 21366
rect 13697 21298 13817 21332
rect 13697 21264 13739 21298
rect 13773 21264 13817 21298
rect 13697 21230 13817 21264
rect 13697 21196 13739 21230
rect 13773 21196 13817 21230
rect 13697 21162 13817 21196
rect 13697 21128 13739 21162
rect 13773 21128 13817 21162
rect 13697 21094 13817 21128
rect 13697 21060 13739 21094
rect 13773 21060 13817 21094
rect 13697 21026 13817 21060
rect 13697 20992 13739 21026
rect 13773 20992 13817 21026
rect 13697 20958 13817 20992
rect 13697 20924 13739 20958
rect 13773 20924 13817 20958
rect 13697 20890 13817 20924
rect 13697 20856 13739 20890
rect 13773 20856 13817 20890
rect 13697 20822 13817 20856
rect 13697 20788 13739 20822
rect 13773 20788 13817 20822
rect 13697 20754 13817 20788
rect 13697 20720 13739 20754
rect 13773 20720 13817 20754
rect 13697 20686 13817 20720
rect 13697 20652 13739 20686
rect 13773 20652 13817 20686
rect 13697 20618 13817 20652
rect 13697 20584 13739 20618
rect 13773 20584 13817 20618
rect 13697 20550 13817 20584
rect 13697 20516 13739 20550
rect 13773 20516 13817 20550
rect 13697 20482 13817 20516
rect 13697 20448 13739 20482
rect 13773 20448 13817 20482
rect 13697 20414 13817 20448
rect 13697 20380 13739 20414
rect 13773 20380 13817 20414
rect 13697 20346 13817 20380
rect 13697 20312 13739 20346
rect 13773 20312 13817 20346
rect 13697 20278 13817 20312
rect 13697 20244 13739 20278
rect 13773 20244 13817 20278
rect 13697 20210 13817 20244
rect 13697 20176 13739 20210
rect 13773 20176 13817 20210
rect 13697 20142 13817 20176
rect 13697 20108 13739 20142
rect 13773 20108 13817 20142
rect 13697 20074 13817 20108
rect 13697 20040 13739 20074
rect 13773 20040 13817 20074
rect 13697 20006 13817 20040
rect 13697 19972 13739 20006
rect 13773 19972 13817 20006
rect 13697 19938 13817 19972
rect 13697 19904 13739 19938
rect 13773 19904 13817 19938
rect 13697 19870 13817 19904
rect 13697 19836 13739 19870
rect 13773 19836 13817 19870
rect 13697 19802 13817 19836
rect 13697 19768 13739 19802
rect 13773 19768 13817 19802
rect 13697 19734 13817 19768
rect 13697 19700 13739 19734
rect 13773 19700 13817 19734
rect 13697 19666 13817 19700
rect 13697 19632 13739 19666
rect 13773 19632 13817 19666
rect 13697 19598 13817 19632
rect 13697 19564 13739 19598
rect 13773 19564 13817 19598
rect 13697 19530 13817 19564
rect 13697 19496 13739 19530
rect 13773 19496 13817 19530
rect 13697 19462 13817 19496
rect 13697 19428 13739 19462
rect 13773 19428 13817 19462
rect 13697 19394 13817 19428
rect 13697 19360 13739 19394
rect 13773 19360 13817 19394
rect 13697 19326 13817 19360
rect 13697 19292 13739 19326
rect 13773 19292 13817 19326
rect 13697 19258 13817 19292
rect 13697 19224 13739 19258
rect 13773 19224 13817 19258
rect 13697 19190 13817 19224
rect 13697 19156 13739 19190
rect 13773 19156 13817 19190
rect 13697 19122 13817 19156
rect 13697 19088 13739 19122
rect 13773 19088 13817 19122
rect 13697 19054 13817 19088
rect 13697 19020 13739 19054
rect 13773 19020 13817 19054
rect 13697 18986 13817 19020
rect 13697 18952 13739 18986
rect 13773 18952 13817 18986
rect 13697 18918 13817 18952
rect 13697 18884 13739 18918
rect 13773 18884 13817 18918
rect 13697 18850 13817 18884
rect 13697 18816 13739 18850
rect 13773 18816 13817 18850
rect 13697 18782 13817 18816
rect 13697 18748 13739 18782
rect 13773 18748 13817 18782
rect 13697 18714 13817 18748
rect 13697 18680 13739 18714
rect 13773 18680 13817 18714
rect 13697 18646 13817 18680
rect 13697 18612 13739 18646
rect 13773 18612 13817 18646
rect 13697 18578 13817 18612
rect 13697 18544 13739 18578
rect 13773 18544 13817 18578
rect 13697 18510 13817 18544
rect 13697 18476 13739 18510
rect 13773 18476 13817 18510
rect 13697 18442 13817 18476
rect 13697 18408 13739 18442
rect 13773 18408 13817 18442
rect 13697 18374 13817 18408
rect 13697 18340 13739 18374
rect 13773 18340 13817 18374
rect 13697 18306 13817 18340
rect 13697 18272 13739 18306
rect 13773 18272 13817 18306
rect 13697 18238 13817 18272
rect 13697 18204 13739 18238
rect 13773 18204 13817 18238
rect 13697 18170 13817 18204
rect 13697 18136 13739 18170
rect 13773 18136 13817 18170
rect 13697 18102 13817 18136
rect 13697 18068 13739 18102
rect 13773 18068 13817 18102
rect 13697 18034 13817 18068
rect 13697 18000 13739 18034
rect 13773 18000 13817 18034
rect 13697 17966 13817 18000
rect 13697 17932 13739 17966
rect 13773 17932 13817 17966
rect 13697 17898 13817 17932
rect 13697 17864 13739 17898
rect 13773 17864 13817 17898
rect 13697 17830 13817 17864
rect 13697 17796 13739 17830
rect 13773 17796 13817 17830
rect 13697 17762 13817 17796
rect 13697 17728 13739 17762
rect 13773 17728 13817 17762
rect 13697 17694 13817 17728
rect 13697 17660 13739 17694
rect 13773 17660 13817 17694
rect 13697 17626 13817 17660
rect 13697 17592 13739 17626
rect 13773 17592 13817 17626
rect 13697 17558 13817 17592
rect 13697 17524 13739 17558
rect 13773 17524 13817 17558
rect 13697 17490 13817 17524
rect 13697 17456 13739 17490
rect 13773 17456 13817 17490
rect 13697 17422 13817 17456
rect 13697 17388 13739 17422
rect 13773 17388 13817 17422
rect 13697 17354 13817 17388
rect 13697 17320 13739 17354
rect 13773 17320 13817 17354
rect 13697 17286 13817 17320
rect 13697 17252 13739 17286
rect 13773 17252 13817 17286
rect 13697 17218 13817 17252
rect 13697 17184 13739 17218
rect 13773 17184 13817 17218
rect 13697 17150 13817 17184
rect 13697 17116 13739 17150
rect 13773 17116 13817 17150
rect 13697 17082 13817 17116
rect 13697 17048 13739 17082
rect 13773 17048 13817 17082
rect 13697 17014 13817 17048
rect 13697 16980 13739 17014
rect 13773 16980 13817 17014
rect 13697 16946 13817 16980
rect 13697 16912 13739 16946
rect 13773 16912 13817 16946
rect 13697 16878 13817 16912
rect 13697 16844 13739 16878
rect 13773 16844 13817 16878
rect 13697 16810 13817 16844
rect 13697 16776 13739 16810
rect 13773 16776 13817 16810
rect 13697 16742 13817 16776
rect 13697 16708 13739 16742
rect 13773 16708 13817 16742
rect 13697 16674 13817 16708
rect 13697 16640 13739 16674
rect 13773 16640 13817 16674
rect 13697 16606 13817 16640
rect 13697 16572 13739 16606
rect 13773 16572 13817 16606
rect 13697 16538 13817 16572
rect 13697 16504 13739 16538
rect 13773 16504 13817 16538
rect 13697 16470 13817 16504
rect 13697 16436 13739 16470
rect 13773 16436 13817 16470
rect 13697 16402 13817 16436
rect 13697 16368 13739 16402
rect 13773 16368 13817 16402
rect 13697 16334 13817 16368
rect 13697 16300 13739 16334
rect 13773 16300 13817 16334
rect 13697 16266 13817 16300
rect 13697 16232 13739 16266
rect 13773 16232 13817 16266
rect 13697 16198 13817 16232
rect 13697 16164 13739 16198
rect 13773 16164 13817 16198
rect 13697 16130 13817 16164
rect 13697 16096 13739 16130
rect 13773 16096 13817 16130
rect 13697 16062 13817 16096
rect 13697 16028 13739 16062
rect 13773 16028 13817 16062
rect 13697 15994 13817 16028
rect 13697 15960 13739 15994
rect 13773 15960 13817 15994
rect 13697 15926 13817 15960
rect 13697 15892 13739 15926
rect 13773 15892 13817 15926
rect 13697 15858 13817 15892
rect 13697 15824 13739 15858
rect 13773 15824 13817 15858
rect 13697 15790 13817 15824
rect 13697 15756 13739 15790
rect 13773 15756 13817 15790
rect 13697 15722 13817 15756
rect 13697 15688 13739 15722
rect 13773 15688 13817 15722
rect 13697 15654 13817 15688
rect 13697 15620 13739 15654
rect 13773 15620 13817 15654
rect 13697 15586 13817 15620
rect 13697 15552 13739 15586
rect 13773 15552 13817 15586
rect 13697 15518 13817 15552
rect 13697 15484 13739 15518
rect 13773 15484 13817 15518
rect 13697 15450 13817 15484
rect 13697 15416 13739 15450
rect 13773 15416 13817 15450
rect 13697 15382 13817 15416
rect 13697 15348 13739 15382
rect 13773 15348 13817 15382
rect 13697 15314 13817 15348
rect 13697 15280 13739 15314
rect 13773 15280 13817 15314
rect 13697 15246 13817 15280
rect 13697 15212 13739 15246
rect 13773 15212 13817 15246
rect 13697 15178 13817 15212
rect 13697 15144 13739 15178
rect 13773 15144 13817 15178
rect 13697 15110 13817 15144
rect 13697 15076 13739 15110
rect 13773 15076 13817 15110
rect 13697 15042 13817 15076
rect 13697 15008 13739 15042
rect 13773 15008 13817 15042
rect 13697 14974 13817 15008
rect 13697 14940 13739 14974
rect 13773 14940 13817 14974
rect 13697 14906 13817 14940
rect 13697 14872 13739 14906
rect 13773 14872 13817 14906
rect 13697 14838 13817 14872
rect 13697 14804 13739 14838
rect 13773 14804 13817 14838
rect 13697 14770 13817 14804
rect 13697 14736 13739 14770
rect 13773 14736 13817 14770
rect 13697 14702 13817 14736
rect 13697 14668 13739 14702
rect 13773 14668 13817 14702
rect 13697 14634 13817 14668
rect 13697 14600 13739 14634
rect 13773 14600 13817 14634
rect 13697 14566 13817 14600
rect 13697 14532 13739 14566
rect 13773 14532 13817 14566
rect 13697 14498 13817 14532
rect 13697 14464 13739 14498
rect 13773 14464 13817 14498
rect 13697 14430 13817 14464
rect 13697 14396 13739 14430
rect 13773 14396 13817 14430
rect 13697 14362 13817 14396
rect 13697 14328 13739 14362
rect 13773 14328 13817 14362
rect 13697 14294 13817 14328
rect 13697 14260 13739 14294
rect 13773 14260 13817 14294
rect 13697 14226 13817 14260
rect 13697 14192 13739 14226
rect 13773 14192 13817 14226
rect 13697 14158 13817 14192
rect 13697 14124 13739 14158
rect 13773 14124 13817 14158
rect 13697 14090 13817 14124
rect 13697 14056 13739 14090
rect 13773 14056 13817 14090
rect 13697 14022 13817 14056
rect 13697 13988 13739 14022
rect 13773 13988 13817 14022
rect 13697 13954 13817 13988
rect 13697 13920 13739 13954
rect 13773 13920 13817 13954
rect 13697 13886 13817 13920
rect 13697 13852 13739 13886
rect 13773 13852 13817 13886
rect 13697 13818 13817 13852
rect 13697 13784 13739 13818
rect 13773 13784 13817 13818
rect 13697 13750 13817 13784
rect 13697 13716 13739 13750
rect 13773 13716 13817 13750
rect 13697 13682 13817 13716
rect 13697 13648 13739 13682
rect 13773 13648 13817 13682
rect 13697 13614 13817 13648
rect 13697 13580 13739 13614
rect 13773 13580 13817 13614
rect 13697 13546 13817 13580
rect 13697 13512 13739 13546
rect 13773 13512 13817 13546
rect 13697 13478 13817 13512
rect 13697 13444 13739 13478
rect 13773 13444 13817 13478
rect 13697 13410 13817 13444
rect 13697 13376 13739 13410
rect 13773 13376 13817 13410
rect 13697 13342 13817 13376
rect 13697 13308 13739 13342
rect 13773 13308 13817 13342
rect 13697 13274 13817 13308
rect 13697 13240 13739 13274
rect 13773 13240 13817 13274
rect 13697 13206 13817 13240
rect 13697 13172 13739 13206
rect 13773 13172 13817 13206
rect 13697 13138 13817 13172
rect 13697 13104 13739 13138
rect 13773 13104 13817 13138
rect 13697 13070 13817 13104
rect 13697 13036 13739 13070
rect 13773 13036 13817 13070
rect 13697 13002 13817 13036
rect 13697 12968 13739 13002
rect 13773 12968 13817 13002
rect 13697 12934 13817 12968
rect 13697 12900 13739 12934
rect 13773 12900 13817 12934
rect 13697 12866 13817 12900
rect 13697 12832 13739 12866
rect 13773 12832 13817 12866
rect 13697 12798 13817 12832
rect 13697 12764 13739 12798
rect 13773 12764 13817 12798
rect 13697 12730 13817 12764
rect 13697 12696 13739 12730
rect 13773 12696 13817 12730
rect 13697 12662 13817 12696
rect 13697 12628 13739 12662
rect 13773 12628 13817 12662
rect 13697 12594 13817 12628
rect 13697 12560 13739 12594
rect 13773 12560 13817 12594
rect 13697 12526 13817 12560
rect 13697 12492 13739 12526
rect 13773 12492 13817 12526
rect 13697 12458 13817 12492
rect 13697 12424 13739 12458
rect 13773 12424 13817 12458
rect 13697 12390 13817 12424
rect 13697 12356 13739 12390
rect 13773 12356 13817 12390
rect 13697 12322 13817 12356
rect 13697 12288 13739 12322
rect 13773 12288 13817 12322
rect 13697 12254 13817 12288
rect 13697 12220 13739 12254
rect 13773 12220 13817 12254
rect 13697 12186 13817 12220
rect 13697 12152 13739 12186
rect 13773 12152 13817 12186
rect 13697 12118 13817 12152
rect 13697 12084 13739 12118
rect 13773 12084 13817 12118
rect 13697 12050 13817 12084
rect 13697 12016 13739 12050
rect 13773 12016 13817 12050
rect 13697 11982 13817 12016
rect 13697 11948 13739 11982
rect 13773 11948 13817 11982
rect 13697 11914 13817 11948
rect 13697 11880 13739 11914
rect 13773 11880 13817 11914
rect 13697 11846 13817 11880
rect 13697 11812 13739 11846
rect 13773 11812 13817 11846
rect 13697 11778 13817 11812
rect 13697 11744 13739 11778
rect 13773 11744 13817 11778
rect 13697 11710 13817 11744
rect 13697 11676 13739 11710
rect 13773 11676 13817 11710
rect 13697 11642 13817 11676
rect 13697 11608 13739 11642
rect 13773 11608 13817 11642
rect 13697 11574 13817 11608
rect 13697 11540 13739 11574
rect 13773 11540 13817 11574
rect 13697 11506 13817 11540
rect 13697 11472 13739 11506
rect 13773 11472 13817 11506
rect 13697 11438 13817 11472
rect 13697 11404 13739 11438
rect 13773 11404 13817 11438
rect 13697 11370 13817 11404
rect 13697 11336 13739 11370
rect 13773 11336 13817 11370
rect 13697 11302 13817 11336
rect 13697 11268 13739 11302
rect 13773 11268 13817 11302
rect 13697 11234 13817 11268
rect 13697 11200 13739 11234
rect 13773 11200 13817 11234
rect 13697 11166 13817 11200
rect 13697 11132 13739 11166
rect 13773 11132 13817 11166
rect 13697 11098 13817 11132
rect 13697 11064 13739 11098
rect 13773 11064 13817 11098
rect 13697 11030 13817 11064
rect 13697 10996 13739 11030
rect 13773 10996 13817 11030
rect 13697 10962 13817 10996
rect 13697 10928 13739 10962
rect 13773 10928 13817 10962
rect 13697 10894 13817 10928
rect 13697 10860 13739 10894
rect 13773 10860 13817 10894
rect 13697 10826 13817 10860
rect 13697 10792 13739 10826
rect 13773 10792 13817 10826
rect 13697 10758 13817 10792
rect 13697 10724 13739 10758
rect 13773 10724 13817 10758
rect 13697 10690 13817 10724
rect 13697 10656 13739 10690
rect 13773 10656 13817 10690
rect 13697 10622 13817 10656
rect 13697 10588 13739 10622
rect 13773 10588 13817 10622
rect 13697 10554 13817 10588
rect 13697 10520 13739 10554
rect 13773 10520 13817 10554
rect 13697 10486 13817 10520
rect 13697 10452 13739 10486
rect 13773 10452 13817 10486
rect 13697 10418 13817 10452
rect 13697 10384 13739 10418
rect 13773 10384 13817 10418
rect 13697 10334 13817 10384
rect 1177 10290 13817 10334
rect 1177 10256 1355 10290
rect 1389 10256 1423 10290
rect 1457 10256 1491 10290
rect 1525 10256 1559 10290
rect 1593 10256 1627 10290
rect 1661 10256 1695 10290
rect 1729 10256 1763 10290
rect 1797 10256 1831 10290
rect 1865 10256 1899 10290
rect 1933 10256 1967 10290
rect 2001 10256 2035 10290
rect 2069 10256 2103 10290
rect 2137 10256 2171 10290
rect 2205 10256 2239 10290
rect 2273 10256 2307 10290
rect 2341 10256 2375 10290
rect 2409 10256 2443 10290
rect 2477 10256 2511 10290
rect 2545 10256 2579 10290
rect 2613 10256 2647 10290
rect 2681 10256 2715 10290
rect 2749 10256 2783 10290
rect 2817 10256 2851 10290
rect 2885 10256 2919 10290
rect 2953 10256 2987 10290
rect 3021 10256 3055 10290
rect 3089 10256 3123 10290
rect 3157 10256 3191 10290
rect 3225 10256 3259 10290
rect 3293 10256 3327 10290
rect 3361 10256 3395 10290
rect 3429 10256 3463 10290
rect 3497 10256 3531 10290
rect 3565 10256 3599 10290
rect 3633 10256 3667 10290
rect 3701 10256 3735 10290
rect 3769 10256 3803 10290
rect 3837 10256 3871 10290
rect 3905 10256 3939 10290
rect 3973 10256 4007 10290
rect 4041 10256 4075 10290
rect 4109 10256 4143 10290
rect 4177 10256 4211 10290
rect 4245 10256 4279 10290
rect 4313 10256 4347 10290
rect 4381 10256 4415 10290
rect 4449 10256 4483 10290
rect 4517 10256 4551 10290
rect 4585 10256 4619 10290
rect 4653 10256 4687 10290
rect 4721 10256 4755 10290
rect 4789 10256 4823 10290
rect 4857 10256 4891 10290
rect 4925 10256 4959 10290
rect 4993 10256 5027 10290
rect 5061 10256 5095 10290
rect 5129 10256 5163 10290
rect 5197 10256 5231 10290
rect 5265 10256 5299 10290
rect 5333 10256 5367 10290
rect 5401 10256 5435 10290
rect 5469 10256 5503 10290
rect 5537 10256 5571 10290
rect 5605 10256 5639 10290
rect 5673 10256 5707 10290
rect 5741 10256 5775 10290
rect 5809 10256 5843 10290
rect 5877 10256 5911 10290
rect 5945 10256 5979 10290
rect 6013 10256 6047 10290
rect 6081 10256 6115 10290
rect 6149 10256 6183 10290
rect 6217 10256 6251 10290
rect 6285 10256 6319 10290
rect 6353 10256 6387 10290
rect 6421 10256 6455 10290
rect 6489 10256 6523 10290
rect 6557 10256 6591 10290
rect 6625 10256 6659 10290
rect 6693 10256 6727 10290
rect 6761 10256 6795 10290
rect 6829 10256 6863 10290
rect 6897 10256 6931 10290
rect 6965 10256 6999 10290
rect 7033 10256 7067 10290
rect 7101 10256 7135 10290
rect 7169 10256 7203 10290
rect 7237 10256 7271 10290
rect 7305 10256 7339 10290
rect 7373 10256 7407 10290
rect 7441 10256 7475 10290
rect 7509 10256 7543 10290
rect 7577 10256 7611 10290
rect 7645 10256 7679 10290
rect 7713 10256 7747 10290
rect 7781 10256 7815 10290
rect 7849 10256 7883 10290
rect 7917 10256 7951 10290
rect 7985 10256 8019 10290
rect 8053 10256 8087 10290
rect 8121 10256 8155 10290
rect 8189 10256 8223 10290
rect 8257 10256 8291 10290
rect 8325 10256 8359 10290
rect 8393 10256 8427 10290
rect 8461 10256 8495 10290
rect 8529 10256 8563 10290
rect 8597 10256 8631 10290
rect 8665 10256 8699 10290
rect 8733 10256 8767 10290
rect 8801 10256 8835 10290
rect 8869 10256 8903 10290
rect 8937 10256 8971 10290
rect 9005 10256 9039 10290
rect 9073 10256 9107 10290
rect 9141 10256 9175 10290
rect 9209 10256 9243 10290
rect 9277 10256 9311 10290
rect 9345 10256 9379 10290
rect 9413 10256 9447 10290
rect 9481 10256 9515 10290
rect 9549 10256 9583 10290
rect 9617 10256 9651 10290
rect 9685 10256 9719 10290
rect 9753 10256 9787 10290
rect 9821 10256 9855 10290
rect 9889 10256 9923 10290
rect 9957 10256 9991 10290
rect 10025 10256 10059 10290
rect 10093 10256 10127 10290
rect 10161 10256 10195 10290
rect 10229 10256 10263 10290
rect 10297 10256 10331 10290
rect 10365 10256 10399 10290
rect 10433 10256 10467 10290
rect 10501 10256 10535 10290
rect 10569 10256 10603 10290
rect 10637 10256 10671 10290
rect 10705 10256 10739 10290
rect 10773 10256 10807 10290
rect 10841 10256 10875 10290
rect 10909 10256 10943 10290
rect 10977 10256 11011 10290
rect 11045 10256 11079 10290
rect 11113 10256 11147 10290
rect 11181 10256 11215 10290
rect 11249 10256 11283 10290
rect 11317 10256 11351 10290
rect 11385 10256 11419 10290
rect 11453 10256 11487 10290
rect 11521 10256 11555 10290
rect 11589 10256 11623 10290
rect 11657 10256 11691 10290
rect 11725 10256 11759 10290
rect 11793 10256 11827 10290
rect 11861 10256 11895 10290
rect 11929 10256 11963 10290
rect 11997 10256 12031 10290
rect 12065 10256 12099 10290
rect 12133 10256 12167 10290
rect 12201 10256 12235 10290
rect 12269 10256 12303 10290
rect 12337 10256 12371 10290
rect 12405 10256 12439 10290
rect 12473 10256 12507 10290
rect 12541 10256 12575 10290
rect 12609 10256 12643 10290
rect 12677 10256 12711 10290
rect 12745 10256 12779 10290
rect 12813 10256 12847 10290
rect 12881 10256 12915 10290
rect 12949 10256 12983 10290
rect 13017 10256 13051 10290
rect 13085 10256 13119 10290
rect 13153 10256 13187 10290
rect 13221 10256 13255 10290
rect 13289 10256 13323 10290
rect 13357 10256 13391 10290
rect 13425 10256 13459 10290
rect 13493 10256 13527 10290
rect 13561 10256 13595 10290
rect 13629 10256 13817 10290
rect 1177 10214 13817 10256
rect 14539 36225 14609 36259
rect 14643 36225 14724 36259
rect 14539 36191 14724 36225
rect 14539 36157 14609 36191
rect 14643 36157 14724 36191
rect 14539 36123 14724 36157
rect 14539 36089 14609 36123
rect 14643 36089 14724 36123
rect 14539 36055 14724 36089
rect 14539 36021 14609 36055
rect 14643 36021 14724 36055
rect 14539 35987 14724 36021
rect 14539 35953 14609 35987
rect 14643 35953 14724 35987
rect 14539 35919 14724 35953
rect 14539 35885 14609 35919
rect 14643 35885 14724 35919
rect 14539 35851 14724 35885
rect 14539 35817 14609 35851
rect 14643 35817 14724 35851
rect 14539 35783 14724 35817
rect 14539 35749 14609 35783
rect 14643 35749 14724 35783
rect 14539 35715 14724 35749
rect 14539 35681 14609 35715
rect 14643 35681 14724 35715
rect 14539 35647 14724 35681
rect 14539 35613 14609 35647
rect 14643 35613 14724 35647
rect 14539 35579 14724 35613
rect 14539 35545 14609 35579
rect 14643 35545 14724 35579
rect 14539 35511 14724 35545
rect 14539 35477 14609 35511
rect 14643 35477 14724 35511
rect 14539 35443 14724 35477
rect 14539 35409 14609 35443
rect 14643 35409 14724 35443
rect 14539 35375 14724 35409
rect 14539 35341 14609 35375
rect 14643 35341 14724 35375
rect 14539 35307 14724 35341
rect 14539 35273 14609 35307
rect 14643 35273 14724 35307
rect 14539 35239 14724 35273
rect 14539 35205 14609 35239
rect 14643 35205 14724 35239
rect 14539 35171 14724 35205
rect 14539 35137 14609 35171
rect 14643 35137 14724 35171
rect 14539 35103 14724 35137
rect 14539 35069 14609 35103
rect 14643 35069 14724 35103
rect 14539 35035 14724 35069
rect 14539 35001 14609 35035
rect 14643 35001 14724 35035
rect 14539 34967 14724 35001
rect 14539 34933 14609 34967
rect 14643 34933 14724 34967
rect 14539 34899 14724 34933
rect 14539 34865 14609 34899
rect 14643 34865 14724 34899
rect 14539 34831 14724 34865
rect 14539 34797 14609 34831
rect 14643 34797 14724 34831
rect 14539 34763 14724 34797
rect 14539 34729 14609 34763
rect 14643 34729 14724 34763
rect 14539 34695 14724 34729
rect 14539 34661 14609 34695
rect 14643 34661 14724 34695
rect 14539 34627 14724 34661
rect 14539 34593 14609 34627
rect 14643 34593 14724 34627
rect 14539 34559 14724 34593
rect 14539 34525 14609 34559
rect 14643 34525 14724 34559
rect 14539 34491 14724 34525
rect 14539 34457 14609 34491
rect 14643 34457 14724 34491
rect 14539 34423 14724 34457
rect 14539 34389 14609 34423
rect 14643 34389 14724 34423
rect 14539 34355 14724 34389
rect 14539 34321 14609 34355
rect 14643 34321 14724 34355
rect 14539 34287 14724 34321
rect 14539 34253 14609 34287
rect 14643 34253 14724 34287
rect 14539 34219 14724 34253
rect 14539 34185 14609 34219
rect 14643 34185 14724 34219
rect 14539 34151 14724 34185
rect 14539 34117 14609 34151
rect 14643 34117 14724 34151
rect 14539 34083 14724 34117
rect 14539 34049 14609 34083
rect 14643 34049 14724 34083
rect 14539 34015 14724 34049
rect 14539 33981 14609 34015
rect 14643 33981 14724 34015
rect 14539 33947 14724 33981
rect 14539 33913 14609 33947
rect 14643 33913 14724 33947
rect 14539 33879 14724 33913
rect 14539 33845 14609 33879
rect 14643 33845 14724 33879
rect 14539 33811 14724 33845
rect 14539 33777 14609 33811
rect 14643 33777 14724 33811
rect 14539 33743 14724 33777
rect 14539 33709 14609 33743
rect 14643 33709 14724 33743
rect 14539 33675 14724 33709
rect 14539 33641 14609 33675
rect 14643 33641 14724 33675
rect 14539 33607 14724 33641
rect 14539 33573 14609 33607
rect 14643 33573 14724 33607
rect 14539 33539 14724 33573
rect 14539 33505 14609 33539
rect 14643 33505 14724 33539
rect 14539 33471 14724 33505
rect 14539 33437 14609 33471
rect 14643 33437 14724 33471
rect 14539 33403 14724 33437
rect 14539 33369 14609 33403
rect 14643 33369 14724 33403
rect 14539 33335 14724 33369
rect 14539 33301 14609 33335
rect 14643 33301 14724 33335
rect 14539 33267 14724 33301
rect 14539 33233 14609 33267
rect 14643 33233 14724 33267
rect 14539 33199 14724 33233
rect 14539 33165 14609 33199
rect 14643 33165 14724 33199
rect 14539 33131 14724 33165
rect 14539 33097 14609 33131
rect 14643 33097 14724 33131
rect 14539 33063 14724 33097
rect 14539 33029 14609 33063
rect 14643 33029 14724 33063
rect 14539 32995 14724 33029
rect 14539 32961 14609 32995
rect 14643 32961 14724 32995
rect 14539 32927 14724 32961
rect 14539 32893 14609 32927
rect 14643 32893 14724 32927
rect 14539 32859 14724 32893
rect 14539 32825 14609 32859
rect 14643 32825 14724 32859
rect 14539 32791 14724 32825
rect 14539 32757 14609 32791
rect 14643 32757 14724 32791
rect 14539 32723 14724 32757
rect 14539 32689 14609 32723
rect 14643 32689 14724 32723
rect 14539 32655 14724 32689
rect 14539 32621 14609 32655
rect 14643 32621 14724 32655
rect 14539 32587 14724 32621
rect 14539 32553 14609 32587
rect 14643 32553 14724 32587
rect 14539 32519 14724 32553
rect 14539 32485 14609 32519
rect 14643 32485 14724 32519
rect 14539 32451 14724 32485
rect 14539 32417 14609 32451
rect 14643 32417 14724 32451
rect 14539 32383 14724 32417
rect 14539 32349 14609 32383
rect 14643 32349 14724 32383
rect 14539 32315 14724 32349
rect 14539 32281 14609 32315
rect 14643 32281 14724 32315
rect 14539 32247 14724 32281
rect 14539 32213 14609 32247
rect 14643 32213 14724 32247
rect 14539 32179 14724 32213
rect 14539 32145 14609 32179
rect 14643 32145 14724 32179
rect 14539 32111 14724 32145
rect 14539 32077 14609 32111
rect 14643 32077 14724 32111
rect 14539 32043 14724 32077
rect 14539 32009 14609 32043
rect 14643 32009 14724 32043
rect 14539 31975 14724 32009
rect 14539 31941 14609 31975
rect 14643 31941 14724 31975
rect 14539 31907 14724 31941
rect 14539 31873 14609 31907
rect 14643 31873 14724 31907
rect 14539 31839 14724 31873
rect 14539 31805 14609 31839
rect 14643 31805 14724 31839
rect 14539 31771 14724 31805
rect 14539 31737 14609 31771
rect 14643 31737 14724 31771
rect 14539 31703 14724 31737
rect 14539 31669 14609 31703
rect 14643 31669 14724 31703
rect 14539 31635 14724 31669
rect 14539 31601 14609 31635
rect 14643 31601 14724 31635
rect 14539 31567 14724 31601
rect 14539 31533 14609 31567
rect 14643 31533 14724 31567
rect 14539 31499 14724 31533
rect 14539 31465 14609 31499
rect 14643 31465 14724 31499
rect 14539 31431 14724 31465
rect 14539 31397 14609 31431
rect 14643 31397 14724 31431
rect 14539 31363 14724 31397
rect 14539 31329 14609 31363
rect 14643 31329 14724 31363
rect 14539 31295 14724 31329
rect 14539 31261 14609 31295
rect 14643 31261 14724 31295
rect 14539 31227 14724 31261
rect 14539 31193 14609 31227
rect 14643 31193 14724 31227
rect 14539 31159 14724 31193
rect 14539 31125 14609 31159
rect 14643 31125 14724 31159
rect 14539 31091 14724 31125
rect 14539 31057 14609 31091
rect 14643 31057 14724 31091
rect 14539 31023 14724 31057
rect 14539 30989 14609 31023
rect 14643 30989 14724 31023
rect 14539 30955 14724 30989
rect 14539 30921 14609 30955
rect 14643 30921 14724 30955
rect 14539 30887 14724 30921
rect 14539 30853 14609 30887
rect 14643 30853 14724 30887
rect 14539 30819 14724 30853
rect 14539 30785 14609 30819
rect 14643 30785 14724 30819
rect 14539 30751 14724 30785
rect 14539 30717 14609 30751
rect 14643 30717 14724 30751
rect 14539 30683 14724 30717
rect 14539 30649 14609 30683
rect 14643 30649 14724 30683
rect 14539 30615 14724 30649
rect 14539 30581 14609 30615
rect 14643 30581 14724 30615
rect 14539 30547 14724 30581
rect 14539 30513 14609 30547
rect 14643 30513 14724 30547
rect 14539 30479 14724 30513
rect 14539 30445 14609 30479
rect 14643 30445 14724 30479
rect 14539 30411 14724 30445
rect 14539 30377 14609 30411
rect 14643 30377 14724 30411
rect 14539 30343 14724 30377
rect 14539 30309 14609 30343
rect 14643 30309 14724 30343
rect 14539 30275 14724 30309
rect 14539 30241 14609 30275
rect 14643 30241 14724 30275
rect 14539 30207 14724 30241
rect 14539 30173 14609 30207
rect 14643 30173 14724 30207
rect 14539 30139 14724 30173
rect 14539 30105 14609 30139
rect 14643 30105 14724 30139
rect 14539 30071 14724 30105
rect 14539 30037 14609 30071
rect 14643 30037 14724 30071
rect 14539 30003 14724 30037
rect 14539 29969 14609 30003
rect 14643 29969 14724 30003
rect 14539 29935 14724 29969
rect 14539 29901 14609 29935
rect 14643 29901 14724 29935
rect 14539 29867 14724 29901
rect 14539 29833 14609 29867
rect 14643 29833 14724 29867
rect 14539 29799 14724 29833
rect 14539 29765 14609 29799
rect 14643 29765 14724 29799
rect 14539 29731 14724 29765
rect 14539 29697 14609 29731
rect 14643 29697 14724 29731
rect 14539 29663 14724 29697
rect 14539 29629 14609 29663
rect 14643 29629 14724 29663
rect 14539 29595 14724 29629
rect 14539 29561 14609 29595
rect 14643 29561 14724 29595
rect 14539 29527 14724 29561
rect 14539 29493 14609 29527
rect 14643 29493 14724 29527
rect 14539 29459 14724 29493
rect 14539 29425 14609 29459
rect 14643 29425 14724 29459
rect 14539 29391 14724 29425
rect 14539 29357 14609 29391
rect 14643 29357 14724 29391
rect 14539 29323 14724 29357
rect 14539 29289 14609 29323
rect 14643 29289 14724 29323
rect 14539 29255 14724 29289
rect 14539 29221 14609 29255
rect 14643 29221 14724 29255
rect 14539 29187 14724 29221
rect 14539 29153 14609 29187
rect 14643 29153 14724 29187
rect 14539 29119 14724 29153
rect 14539 29085 14609 29119
rect 14643 29085 14724 29119
rect 14539 29051 14724 29085
rect 14539 29017 14609 29051
rect 14643 29017 14724 29051
rect 14539 28983 14724 29017
rect 14539 28949 14609 28983
rect 14643 28949 14724 28983
rect 14539 28915 14724 28949
rect 14539 28881 14609 28915
rect 14643 28881 14724 28915
rect 14539 28847 14724 28881
rect 14539 28813 14609 28847
rect 14643 28813 14724 28847
rect 14539 28779 14724 28813
rect 14539 28745 14609 28779
rect 14643 28745 14724 28779
rect 14539 28711 14724 28745
rect 14539 28677 14609 28711
rect 14643 28677 14724 28711
rect 14539 28643 14724 28677
rect 14539 28609 14609 28643
rect 14643 28609 14724 28643
rect 14539 28575 14724 28609
rect 14539 28541 14609 28575
rect 14643 28541 14724 28575
rect 14539 28507 14724 28541
rect 14539 28473 14609 28507
rect 14643 28473 14724 28507
rect 14539 28439 14724 28473
rect 14539 28405 14609 28439
rect 14643 28405 14724 28439
rect 14539 28371 14724 28405
rect 14539 28337 14609 28371
rect 14643 28337 14724 28371
rect 14539 28303 14724 28337
rect 14539 28269 14609 28303
rect 14643 28269 14724 28303
rect 14539 28235 14724 28269
rect 14539 28201 14609 28235
rect 14643 28201 14724 28235
rect 14539 28167 14724 28201
rect 14539 28133 14609 28167
rect 14643 28133 14724 28167
rect 14539 28099 14724 28133
rect 14539 28065 14609 28099
rect 14643 28065 14724 28099
rect 14539 28031 14724 28065
rect 14539 27997 14609 28031
rect 14643 27997 14724 28031
rect 14539 27963 14724 27997
rect 14539 27929 14609 27963
rect 14643 27929 14724 27963
rect 14539 27895 14724 27929
rect 14539 27861 14609 27895
rect 14643 27861 14724 27895
rect 14539 27827 14724 27861
rect 14539 27793 14609 27827
rect 14643 27793 14724 27827
rect 14539 27759 14724 27793
rect 14539 27725 14609 27759
rect 14643 27725 14724 27759
rect 14539 27691 14724 27725
rect 14539 27657 14609 27691
rect 14643 27657 14724 27691
rect 14539 27623 14724 27657
rect 14539 27589 14609 27623
rect 14643 27589 14724 27623
rect 14539 27555 14724 27589
rect 14539 27521 14609 27555
rect 14643 27521 14724 27555
rect 14539 27487 14724 27521
rect 14539 27453 14609 27487
rect 14643 27453 14724 27487
rect 14539 27419 14724 27453
rect 14539 27385 14609 27419
rect 14643 27385 14724 27419
rect 14539 27351 14724 27385
rect 14539 27317 14609 27351
rect 14643 27317 14724 27351
rect 14539 27283 14724 27317
rect 14539 27249 14609 27283
rect 14643 27249 14724 27283
rect 14539 27215 14724 27249
rect 14539 27181 14609 27215
rect 14643 27181 14724 27215
rect 14539 27147 14724 27181
rect 14539 27113 14609 27147
rect 14643 27113 14724 27147
rect 14539 27079 14724 27113
rect 14539 27045 14609 27079
rect 14643 27045 14724 27079
rect 14539 27011 14724 27045
rect 14539 26977 14609 27011
rect 14643 26977 14724 27011
rect 14539 26943 14724 26977
rect 14539 26909 14609 26943
rect 14643 26909 14724 26943
rect 14539 26875 14724 26909
rect 14539 26841 14609 26875
rect 14643 26841 14724 26875
rect 14539 26807 14724 26841
rect 14539 26773 14609 26807
rect 14643 26773 14724 26807
rect 14539 26739 14724 26773
rect 14539 26705 14609 26739
rect 14643 26705 14724 26739
rect 14539 26671 14724 26705
rect 14539 26637 14609 26671
rect 14643 26637 14724 26671
rect 14539 26603 14724 26637
rect 14539 26569 14609 26603
rect 14643 26569 14724 26603
rect 14539 26535 14724 26569
rect 14539 26501 14609 26535
rect 14643 26501 14724 26535
rect 14539 26467 14724 26501
rect 14539 26433 14609 26467
rect 14643 26433 14724 26467
rect 14539 26399 14724 26433
rect 14539 26365 14609 26399
rect 14643 26365 14724 26399
rect 14539 26331 14724 26365
rect 14539 26297 14609 26331
rect 14643 26297 14724 26331
rect 14539 26263 14724 26297
rect 14539 26229 14609 26263
rect 14643 26229 14724 26263
rect 14539 26195 14724 26229
rect 14539 26161 14609 26195
rect 14643 26161 14724 26195
rect 14539 26127 14724 26161
rect 14539 26093 14609 26127
rect 14643 26093 14724 26127
rect 14539 26059 14724 26093
rect 14539 26025 14609 26059
rect 14643 26025 14724 26059
rect 14539 25991 14724 26025
rect 14539 25957 14609 25991
rect 14643 25957 14724 25991
rect 14539 25923 14724 25957
rect 14539 25889 14609 25923
rect 14643 25889 14724 25923
rect 14539 25855 14724 25889
rect 14539 25821 14609 25855
rect 14643 25821 14724 25855
rect 14539 25787 14724 25821
rect 14539 25753 14609 25787
rect 14643 25753 14724 25787
rect 14539 25719 14724 25753
rect 14539 25685 14609 25719
rect 14643 25685 14724 25719
rect 14539 25651 14724 25685
rect 14539 25617 14609 25651
rect 14643 25617 14724 25651
rect 14539 25583 14724 25617
rect 14539 25549 14609 25583
rect 14643 25549 14724 25583
rect 14539 25515 14724 25549
rect 14539 25481 14609 25515
rect 14643 25481 14724 25515
rect 14539 25447 14724 25481
rect 14539 25413 14609 25447
rect 14643 25413 14724 25447
rect 14539 25379 14724 25413
rect 14539 25345 14609 25379
rect 14643 25345 14724 25379
rect 14539 25311 14724 25345
rect 14539 25277 14609 25311
rect 14643 25277 14724 25311
rect 14539 25243 14724 25277
rect 14539 25209 14609 25243
rect 14643 25209 14724 25243
rect 14539 25175 14724 25209
rect 14539 25141 14609 25175
rect 14643 25141 14724 25175
rect 14539 25107 14724 25141
rect 14539 25073 14609 25107
rect 14643 25073 14724 25107
rect 14539 25039 14724 25073
rect 14539 25005 14609 25039
rect 14643 25005 14724 25039
rect 14539 24971 14724 25005
rect 14539 24937 14609 24971
rect 14643 24937 14724 24971
rect 14539 24903 14724 24937
rect 14539 24869 14609 24903
rect 14643 24869 14724 24903
rect 14539 24835 14724 24869
rect 14539 24801 14609 24835
rect 14643 24801 14724 24835
rect 14539 24767 14724 24801
rect 14539 24733 14609 24767
rect 14643 24733 14724 24767
rect 14539 24699 14724 24733
rect 14539 24665 14609 24699
rect 14643 24665 14724 24699
rect 14539 24631 14724 24665
rect 14539 24597 14609 24631
rect 14643 24597 14724 24631
rect 14539 24563 14724 24597
rect 14539 24529 14609 24563
rect 14643 24529 14724 24563
rect 14539 24495 14724 24529
rect 14539 24461 14609 24495
rect 14643 24461 14724 24495
rect 14539 24427 14724 24461
rect 14539 24393 14609 24427
rect 14643 24393 14724 24427
rect 14539 24359 14724 24393
rect 14539 24325 14609 24359
rect 14643 24325 14724 24359
rect 14539 24291 14724 24325
rect 14539 24257 14609 24291
rect 14643 24257 14724 24291
rect 14539 24223 14724 24257
rect 14539 24189 14609 24223
rect 14643 24189 14724 24223
rect 14539 24155 14724 24189
rect 14539 24121 14609 24155
rect 14643 24121 14724 24155
rect 14539 24087 14724 24121
rect 14539 24053 14609 24087
rect 14643 24053 14724 24087
rect 14539 24019 14724 24053
rect 14539 23985 14609 24019
rect 14643 23985 14724 24019
rect 14539 23951 14724 23985
rect 14539 23917 14609 23951
rect 14643 23917 14724 23951
rect 14539 23883 14724 23917
rect 14539 23849 14609 23883
rect 14643 23849 14724 23883
rect 14539 23815 14724 23849
rect 14539 23781 14609 23815
rect 14643 23781 14724 23815
rect 14539 23747 14724 23781
rect 14539 23713 14609 23747
rect 14643 23713 14724 23747
rect 14539 23679 14724 23713
rect 14539 23645 14609 23679
rect 14643 23645 14724 23679
rect 14539 23611 14724 23645
rect 14539 23577 14609 23611
rect 14643 23577 14724 23611
rect 14539 23543 14724 23577
rect 14539 23509 14609 23543
rect 14643 23509 14724 23543
rect 14539 23475 14724 23509
rect 14539 23441 14609 23475
rect 14643 23441 14724 23475
rect 14539 23407 14724 23441
rect 14539 23373 14609 23407
rect 14643 23373 14724 23407
rect 14539 23339 14724 23373
rect 14539 23305 14609 23339
rect 14643 23305 14724 23339
rect 14539 23271 14724 23305
rect 14539 23237 14609 23271
rect 14643 23237 14724 23271
rect 14539 23203 14724 23237
rect 14539 23169 14609 23203
rect 14643 23169 14724 23203
rect 14539 23135 14724 23169
rect 14539 23101 14609 23135
rect 14643 23101 14724 23135
rect 14539 23067 14724 23101
rect 14539 23033 14609 23067
rect 14643 23033 14724 23067
rect 14539 22999 14724 23033
rect 14539 22965 14609 22999
rect 14643 22965 14724 22999
rect 14539 22931 14724 22965
rect 14539 22897 14609 22931
rect 14643 22897 14724 22931
rect 14539 22863 14724 22897
rect 14539 22829 14609 22863
rect 14643 22829 14724 22863
rect 14539 22795 14724 22829
rect 14539 22761 14609 22795
rect 14643 22761 14724 22795
rect 14539 22727 14724 22761
rect 14539 22693 14609 22727
rect 14643 22693 14724 22727
rect 14539 22659 14724 22693
rect 14539 22625 14609 22659
rect 14643 22625 14724 22659
rect 14539 22591 14724 22625
rect 14539 22557 14609 22591
rect 14643 22557 14724 22591
rect 14539 22523 14724 22557
rect 14539 22489 14609 22523
rect 14643 22489 14724 22523
rect 14539 22455 14724 22489
rect 14539 22421 14609 22455
rect 14643 22421 14724 22455
rect 14539 22387 14724 22421
rect 14539 22353 14609 22387
rect 14643 22353 14724 22387
rect 14539 22319 14724 22353
rect 14539 22285 14609 22319
rect 14643 22285 14724 22319
rect 14539 22251 14724 22285
rect 14539 22217 14609 22251
rect 14643 22217 14724 22251
rect 14539 22183 14724 22217
rect 14539 22149 14609 22183
rect 14643 22149 14724 22183
rect 14539 22115 14724 22149
rect 14539 22081 14609 22115
rect 14643 22081 14724 22115
rect 14539 22047 14724 22081
rect 14539 22013 14609 22047
rect 14643 22013 14724 22047
rect 14539 21979 14724 22013
rect 14539 21945 14609 21979
rect 14643 21945 14724 21979
rect 14539 21911 14724 21945
rect 14539 21877 14609 21911
rect 14643 21877 14724 21911
rect 14539 21843 14724 21877
rect 14539 21809 14609 21843
rect 14643 21809 14724 21843
rect 14539 21775 14724 21809
rect 14539 21741 14609 21775
rect 14643 21741 14724 21775
rect 14539 21707 14724 21741
rect 14539 21673 14609 21707
rect 14643 21673 14724 21707
rect 14539 21639 14724 21673
rect 14539 21605 14609 21639
rect 14643 21605 14724 21639
rect 14539 21571 14724 21605
rect 14539 21537 14609 21571
rect 14643 21537 14724 21571
rect 14539 21503 14724 21537
rect 14539 21469 14609 21503
rect 14643 21469 14724 21503
rect 14539 21435 14724 21469
rect 14539 21401 14609 21435
rect 14643 21401 14724 21435
rect 14539 21367 14724 21401
rect 14539 21333 14609 21367
rect 14643 21333 14724 21367
rect 14539 21299 14724 21333
rect 14539 21265 14609 21299
rect 14643 21265 14724 21299
rect 14539 21231 14724 21265
rect 14539 21197 14609 21231
rect 14643 21197 14724 21231
rect 14539 21163 14724 21197
rect 14539 21129 14609 21163
rect 14643 21129 14724 21163
rect 14539 21095 14724 21129
rect 14539 21061 14609 21095
rect 14643 21061 14724 21095
rect 14539 21027 14724 21061
rect 14539 20993 14609 21027
rect 14643 20993 14724 21027
rect 14539 20959 14724 20993
rect 14539 20925 14609 20959
rect 14643 20925 14724 20959
rect 14539 20891 14724 20925
rect 14539 20857 14609 20891
rect 14643 20857 14724 20891
rect 14539 20823 14724 20857
rect 14539 20789 14609 20823
rect 14643 20789 14724 20823
rect 14539 20755 14724 20789
rect 14539 20721 14609 20755
rect 14643 20721 14724 20755
rect 14539 20687 14724 20721
rect 14539 20653 14609 20687
rect 14643 20653 14724 20687
rect 14539 20619 14724 20653
rect 14539 20585 14609 20619
rect 14643 20585 14724 20619
rect 14539 20551 14724 20585
rect 14539 20517 14609 20551
rect 14643 20517 14724 20551
rect 14539 20483 14724 20517
rect 14539 20449 14609 20483
rect 14643 20449 14724 20483
rect 14539 20415 14724 20449
rect 14539 20381 14609 20415
rect 14643 20381 14724 20415
rect 14539 20347 14724 20381
rect 14539 20313 14609 20347
rect 14643 20313 14724 20347
rect 14539 20279 14724 20313
rect 14539 20245 14609 20279
rect 14643 20245 14724 20279
rect 14539 20211 14724 20245
rect 14539 20177 14609 20211
rect 14643 20177 14724 20211
rect 14539 20143 14724 20177
rect 14539 20109 14609 20143
rect 14643 20109 14724 20143
rect 14539 20075 14724 20109
rect 14539 20041 14609 20075
rect 14643 20041 14724 20075
rect 14539 20007 14724 20041
rect 14539 19973 14609 20007
rect 14643 19973 14724 20007
rect 14539 19939 14724 19973
rect 14539 19905 14609 19939
rect 14643 19905 14724 19939
rect 14539 19871 14724 19905
rect 14539 19837 14609 19871
rect 14643 19837 14724 19871
rect 14539 19803 14724 19837
rect 14539 19769 14609 19803
rect 14643 19769 14724 19803
rect 14539 19735 14724 19769
rect 14539 19701 14609 19735
rect 14643 19701 14724 19735
rect 14539 19667 14724 19701
rect 14539 19633 14609 19667
rect 14643 19633 14724 19667
rect 14539 19599 14724 19633
rect 14539 19565 14609 19599
rect 14643 19565 14724 19599
rect 14539 19531 14724 19565
rect 14539 19497 14609 19531
rect 14643 19497 14724 19531
rect 14539 19463 14724 19497
rect 14539 19429 14609 19463
rect 14643 19429 14724 19463
rect 14539 19395 14724 19429
rect 14539 19361 14609 19395
rect 14643 19361 14724 19395
rect 14539 19327 14724 19361
rect 14539 19293 14609 19327
rect 14643 19293 14724 19327
rect 14539 19259 14724 19293
rect 14539 19225 14609 19259
rect 14643 19225 14724 19259
rect 14539 19191 14724 19225
rect 14539 19157 14609 19191
rect 14643 19157 14724 19191
rect 14539 19123 14724 19157
rect 14539 19089 14609 19123
rect 14643 19089 14724 19123
rect 14539 19055 14724 19089
rect 14539 19021 14609 19055
rect 14643 19021 14724 19055
rect 14539 18987 14724 19021
rect 14539 18953 14609 18987
rect 14643 18953 14724 18987
rect 14539 18919 14724 18953
rect 14539 18885 14609 18919
rect 14643 18885 14724 18919
rect 14539 18851 14724 18885
rect 14539 18817 14609 18851
rect 14643 18817 14724 18851
rect 14539 18783 14724 18817
rect 14539 18749 14609 18783
rect 14643 18749 14724 18783
rect 14539 18715 14724 18749
rect 14539 18681 14609 18715
rect 14643 18681 14724 18715
rect 14539 18647 14724 18681
rect 14539 18613 14609 18647
rect 14643 18613 14724 18647
rect 14539 18579 14724 18613
rect 14539 18545 14609 18579
rect 14643 18545 14724 18579
rect 14539 18511 14724 18545
rect 14539 18477 14609 18511
rect 14643 18477 14724 18511
rect 14539 18443 14724 18477
rect 14539 18409 14609 18443
rect 14643 18409 14724 18443
rect 14539 18375 14724 18409
rect 14539 18341 14609 18375
rect 14643 18341 14724 18375
rect 14539 18307 14724 18341
rect 14539 18273 14609 18307
rect 14643 18273 14724 18307
rect 14539 18239 14724 18273
rect 14539 18205 14609 18239
rect 14643 18205 14724 18239
rect 14539 18171 14724 18205
rect 14539 18137 14609 18171
rect 14643 18137 14724 18171
rect 14539 18103 14724 18137
rect 14539 18069 14609 18103
rect 14643 18069 14724 18103
rect 14539 18035 14724 18069
rect 14539 18001 14609 18035
rect 14643 18001 14724 18035
rect 14539 17967 14724 18001
rect 14539 17933 14609 17967
rect 14643 17933 14724 17967
rect 14539 17899 14724 17933
rect 14539 17865 14609 17899
rect 14643 17865 14724 17899
rect 14539 17831 14724 17865
rect 14539 17797 14609 17831
rect 14643 17797 14724 17831
rect 14539 17763 14724 17797
rect 14539 17729 14609 17763
rect 14643 17729 14724 17763
rect 14539 17695 14724 17729
rect 14539 17661 14609 17695
rect 14643 17661 14724 17695
rect 14539 17627 14724 17661
rect 14539 17593 14609 17627
rect 14643 17593 14724 17627
rect 14539 17559 14724 17593
rect 14539 17525 14609 17559
rect 14643 17525 14724 17559
rect 14539 17491 14724 17525
rect 14539 17457 14609 17491
rect 14643 17457 14724 17491
rect 14539 17423 14724 17457
rect 14539 17389 14609 17423
rect 14643 17389 14724 17423
rect 14539 17355 14724 17389
rect 14539 17321 14609 17355
rect 14643 17321 14724 17355
rect 14539 17287 14724 17321
rect 14539 17253 14609 17287
rect 14643 17253 14724 17287
rect 14539 17219 14724 17253
rect 14539 17185 14609 17219
rect 14643 17185 14724 17219
rect 14539 17151 14724 17185
rect 14539 17117 14609 17151
rect 14643 17117 14724 17151
rect 14539 17083 14724 17117
rect 14539 17049 14609 17083
rect 14643 17049 14724 17083
rect 14539 17015 14724 17049
rect 14539 16981 14609 17015
rect 14643 16981 14724 17015
rect 14539 16947 14724 16981
rect 14539 16913 14609 16947
rect 14643 16913 14724 16947
rect 14539 16879 14724 16913
rect 14539 16845 14609 16879
rect 14643 16845 14724 16879
rect 14539 16811 14724 16845
rect 14539 16777 14609 16811
rect 14643 16777 14724 16811
rect 14539 16743 14724 16777
rect 14539 16709 14609 16743
rect 14643 16709 14724 16743
rect 14539 16675 14724 16709
rect 14539 16641 14609 16675
rect 14643 16641 14724 16675
rect 14539 16607 14724 16641
rect 14539 16573 14609 16607
rect 14643 16573 14724 16607
rect 14539 16539 14724 16573
rect 14539 16505 14609 16539
rect 14643 16505 14724 16539
rect 14539 16471 14724 16505
rect 14539 16437 14609 16471
rect 14643 16437 14724 16471
rect 14539 16403 14724 16437
rect 14539 16369 14609 16403
rect 14643 16369 14724 16403
rect 14539 16335 14724 16369
rect 14539 16301 14609 16335
rect 14643 16301 14724 16335
rect 14539 16267 14724 16301
rect 14539 16233 14609 16267
rect 14643 16233 14724 16267
rect 14539 16199 14724 16233
rect 14539 16165 14609 16199
rect 14643 16165 14724 16199
rect 14539 16131 14724 16165
rect 14539 16097 14609 16131
rect 14643 16097 14724 16131
rect 14539 16063 14724 16097
rect 14539 16029 14609 16063
rect 14643 16029 14724 16063
rect 14539 15995 14724 16029
rect 14539 15961 14609 15995
rect 14643 15961 14724 15995
rect 14539 15927 14724 15961
rect 14539 15893 14609 15927
rect 14643 15893 14724 15927
rect 14539 15859 14724 15893
rect 14539 15825 14609 15859
rect 14643 15825 14724 15859
rect 14539 15791 14724 15825
rect 14539 15757 14609 15791
rect 14643 15757 14724 15791
rect 14539 15723 14724 15757
rect 14539 15689 14609 15723
rect 14643 15689 14724 15723
rect 14539 15655 14724 15689
rect 14539 15621 14609 15655
rect 14643 15621 14724 15655
rect 14539 15587 14724 15621
rect 14539 15553 14609 15587
rect 14643 15553 14724 15587
rect 14539 15519 14724 15553
rect 14539 15485 14609 15519
rect 14643 15485 14724 15519
rect 14539 15451 14724 15485
rect 14539 15417 14609 15451
rect 14643 15417 14724 15451
rect 14539 15383 14724 15417
rect 14539 15349 14609 15383
rect 14643 15349 14724 15383
rect 14539 15315 14724 15349
rect 14539 15281 14609 15315
rect 14643 15281 14724 15315
rect 14539 15247 14724 15281
rect 14539 15213 14609 15247
rect 14643 15213 14724 15247
rect 14539 15179 14724 15213
rect 14539 15145 14609 15179
rect 14643 15145 14724 15179
rect 14539 15111 14724 15145
rect 14539 15077 14609 15111
rect 14643 15077 14724 15111
rect 14539 15043 14724 15077
rect 14539 15009 14609 15043
rect 14643 15009 14724 15043
rect 14539 14975 14724 15009
rect 14539 14941 14609 14975
rect 14643 14941 14724 14975
rect 14539 14907 14724 14941
rect 14539 14873 14609 14907
rect 14643 14873 14724 14907
rect 14539 14839 14724 14873
rect 14539 14805 14609 14839
rect 14643 14805 14724 14839
rect 14539 14771 14724 14805
rect 14539 14737 14609 14771
rect 14643 14737 14724 14771
rect 14539 14703 14724 14737
rect 14539 14669 14609 14703
rect 14643 14669 14724 14703
rect 14539 14635 14724 14669
rect 14539 14601 14609 14635
rect 14643 14601 14724 14635
rect 14539 14567 14724 14601
rect 14539 14533 14609 14567
rect 14643 14533 14724 14567
rect 14539 14499 14724 14533
rect 14539 14465 14609 14499
rect 14643 14465 14724 14499
rect 14539 14431 14724 14465
rect 14539 14397 14609 14431
rect 14643 14397 14724 14431
rect 14539 14363 14724 14397
rect 14539 14329 14609 14363
rect 14643 14329 14724 14363
rect 14539 14295 14724 14329
rect 14539 14261 14609 14295
rect 14643 14261 14724 14295
rect 14539 14227 14724 14261
rect 14539 14193 14609 14227
rect 14643 14193 14724 14227
rect 14539 14159 14724 14193
rect 14539 14125 14609 14159
rect 14643 14125 14724 14159
rect 14539 14091 14724 14125
rect 14539 14057 14609 14091
rect 14643 14057 14724 14091
rect 14539 14023 14724 14057
rect 14539 13989 14609 14023
rect 14643 13989 14724 14023
rect 14539 13955 14724 13989
rect 14539 13921 14609 13955
rect 14643 13921 14724 13955
rect 14539 13887 14724 13921
rect 14539 13853 14609 13887
rect 14643 13853 14724 13887
rect 14539 13819 14724 13853
rect 14539 13785 14609 13819
rect 14643 13785 14724 13819
rect 14539 13751 14724 13785
rect 14539 13717 14609 13751
rect 14643 13717 14724 13751
rect 14539 13683 14724 13717
rect 14539 13649 14609 13683
rect 14643 13649 14724 13683
rect 14539 13615 14724 13649
rect 14539 13581 14609 13615
rect 14643 13581 14724 13615
rect 14539 13547 14724 13581
rect 14539 13513 14609 13547
rect 14643 13513 14724 13547
rect 14539 13479 14724 13513
rect 14539 13445 14609 13479
rect 14643 13445 14724 13479
rect 14539 13411 14724 13445
rect 14539 13377 14609 13411
rect 14643 13377 14724 13411
rect 14539 13343 14724 13377
rect 14539 13309 14609 13343
rect 14643 13309 14724 13343
rect 14539 13275 14724 13309
rect 14539 13241 14609 13275
rect 14643 13241 14724 13275
rect 14539 13207 14724 13241
rect 14539 13173 14609 13207
rect 14643 13173 14724 13207
rect 14539 13139 14724 13173
rect 14539 13105 14609 13139
rect 14643 13105 14724 13139
rect 14539 13071 14724 13105
rect 14539 13037 14609 13071
rect 14643 13037 14724 13071
rect 14539 13003 14724 13037
rect 14539 12969 14609 13003
rect 14643 12969 14724 13003
rect 14539 12935 14724 12969
rect 14539 12901 14609 12935
rect 14643 12901 14724 12935
rect 14539 12867 14724 12901
rect 14539 12833 14609 12867
rect 14643 12833 14724 12867
rect 14539 12799 14724 12833
rect 14539 12765 14609 12799
rect 14643 12765 14724 12799
rect 14539 12731 14724 12765
rect 14539 12697 14609 12731
rect 14643 12697 14724 12731
rect 14539 12663 14724 12697
rect 14539 12629 14609 12663
rect 14643 12629 14724 12663
rect 14539 12595 14724 12629
rect 14539 12561 14609 12595
rect 14643 12561 14724 12595
rect 14539 12527 14724 12561
rect 14539 12493 14609 12527
rect 14643 12493 14724 12527
rect 14539 12459 14724 12493
rect 14539 12425 14609 12459
rect 14643 12425 14724 12459
rect 14539 12391 14724 12425
rect 14539 12357 14609 12391
rect 14643 12357 14724 12391
rect 14539 12323 14724 12357
rect 14539 12289 14609 12323
rect 14643 12289 14724 12323
rect 14539 12255 14724 12289
rect 14539 12221 14609 12255
rect 14643 12221 14724 12255
rect 14539 12187 14724 12221
rect 14539 12153 14609 12187
rect 14643 12153 14724 12187
rect 14539 12119 14724 12153
rect 14539 12085 14609 12119
rect 14643 12085 14724 12119
rect 14539 12051 14724 12085
rect 14539 12017 14609 12051
rect 14643 12017 14724 12051
rect 14539 11983 14724 12017
rect 14539 11949 14609 11983
rect 14643 11949 14724 11983
rect 14539 11915 14724 11949
rect 14539 11881 14609 11915
rect 14643 11881 14724 11915
rect 14539 11847 14724 11881
rect 14539 11813 14609 11847
rect 14643 11813 14724 11847
rect 14539 11779 14724 11813
rect 14539 11745 14609 11779
rect 14643 11745 14724 11779
rect 14539 11711 14724 11745
rect 14539 11677 14609 11711
rect 14643 11677 14724 11711
rect 14539 11643 14724 11677
rect 14539 11609 14609 11643
rect 14643 11609 14724 11643
rect 14539 11575 14724 11609
rect 14539 11541 14609 11575
rect 14643 11541 14724 11575
rect 14539 11507 14724 11541
rect 14539 11473 14609 11507
rect 14643 11473 14724 11507
rect 14539 11439 14724 11473
rect 14539 11405 14609 11439
rect 14643 11405 14724 11439
rect 14539 11371 14724 11405
rect 14539 11337 14609 11371
rect 14643 11337 14724 11371
rect 14539 11303 14724 11337
rect 14539 11269 14609 11303
rect 14643 11269 14724 11303
rect 14539 11235 14724 11269
rect 14539 11201 14609 11235
rect 14643 11201 14724 11235
rect 14539 11167 14724 11201
rect 14539 11133 14609 11167
rect 14643 11133 14724 11167
rect 14539 11099 14724 11133
rect 14539 11065 14609 11099
rect 14643 11065 14724 11099
rect 14539 11031 14724 11065
rect 14539 10997 14609 11031
rect 14643 10997 14724 11031
rect 14539 10963 14724 10997
rect 14539 10929 14609 10963
rect 14643 10929 14724 10963
rect 14539 10895 14724 10929
rect 14539 10861 14609 10895
rect 14643 10861 14724 10895
rect 14539 10827 14724 10861
rect 14539 10793 14609 10827
rect 14643 10793 14724 10827
rect 14539 10759 14724 10793
rect 14539 10725 14609 10759
rect 14643 10725 14724 10759
rect 14539 10691 14724 10725
rect 14539 10657 14609 10691
rect 14643 10657 14724 10691
rect 14539 10623 14724 10657
rect 14539 10589 14609 10623
rect 14643 10589 14724 10623
rect 14539 10555 14724 10589
rect 14539 10521 14609 10555
rect 14643 10521 14724 10555
rect 14539 10487 14724 10521
rect 14539 10453 14609 10487
rect 14643 10453 14724 10487
rect 14539 10419 14724 10453
rect 14539 10385 14609 10419
rect 14643 10385 14724 10419
rect 14539 10351 14724 10385
rect 14539 10317 14609 10351
rect 14643 10317 14724 10351
rect 14539 10283 14724 10317
rect 14539 10249 14609 10283
rect 14643 10249 14724 10283
rect 14539 10215 14724 10249
rect 14539 10181 14609 10215
rect 14643 10181 14724 10215
rect 14539 10147 14724 10181
rect 14539 10113 14609 10147
rect 14643 10113 14724 10147
rect 14539 10079 14724 10113
rect 14539 10045 14609 10079
rect 14643 10045 14724 10079
rect 14539 10011 14724 10045
rect 14539 9977 14609 10011
rect 14643 9977 14724 10011
rect 14539 9943 14724 9977
rect 14539 9909 14609 9943
rect 14643 9909 14724 9943
rect 14539 9875 14724 9909
rect 14539 9841 14609 9875
rect 14643 9841 14724 9875
rect 14539 9807 14724 9841
rect 14539 9773 14609 9807
rect 14643 9773 14724 9807
rect 14539 9739 14724 9773
rect 14539 9705 14609 9739
rect 14643 9705 14724 9739
rect 245 9645 322 9679
rect 356 9645 430 9679
rect 245 9611 430 9645
rect 245 9577 322 9611
rect 356 9577 430 9611
rect 245 9528 430 9577
rect 14539 9671 14724 9705
rect 14539 9637 14609 9671
rect 14643 9637 14724 9671
rect 14539 9603 14724 9637
rect 14539 9569 14609 9603
rect 14643 9569 14724 9603
rect 14539 9528 14724 9569
rect 245 9454 14724 9528
rect 245 9420 510 9454
rect 544 9420 578 9454
rect 612 9420 646 9454
rect 680 9420 714 9454
rect 748 9420 782 9454
rect 816 9420 850 9454
rect 884 9420 918 9454
rect 952 9420 986 9454
rect 1020 9420 1054 9454
rect 1088 9420 1122 9454
rect 1156 9420 1190 9454
rect 1224 9420 1258 9454
rect 1292 9420 1326 9454
rect 1360 9420 1394 9454
rect 1428 9420 1462 9454
rect 1496 9420 1530 9454
rect 1564 9420 1598 9454
rect 1632 9420 1666 9454
rect 1700 9420 1734 9454
rect 1768 9420 1802 9454
rect 1836 9420 1870 9454
rect 1904 9420 1938 9454
rect 1972 9420 2006 9454
rect 2040 9420 2074 9454
rect 2108 9420 2142 9454
rect 2176 9420 2210 9454
rect 2244 9420 2278 9454
rect 2312 9420 2346 9454
rect 2380 9420 2414 9454
rect 2448 9420 2482 9454
rect 2516 9420 2550 9454
rect 2584 9420 2618 9454
rect 2652 9420 2686 9454
rect 2720 9420 2754 9454
rect 2788 9420 2822 9454
rect 2856 9420 2890 9454
rect 2924 9420 2958 9454
rect 2992 9420 3026 9454
rect 3060 9420 3094 9454
rect 3128 9420 3162 9454
rect 3196 9420 3230 9454
rect 3264 9420 3298 9454
rect 3332 9420 3366 9454
rect 3400 9420 3434 9454
rect 3468 9420 3502 9454
rect 3536 9420 3570 9454
rect 3604 9420 3638 9454
rect 3672 9420 3706 9454
rect 3740 9420 3774 9454
rect 3808 9420 3842 9454
rect 3876 9420 3910 9454
rect 3944 9420 3978 9454
rect 4012 9420 4046 9454
rect 4080 9420 4114 9454
rect 4148 9420 4182 9454
rect 4216 9420 4250 9454
rect 4284 9420 4318 9454
rect 4352 9420 4386 9454
rect 4420 9420 4454 9454
rect 4488 9420 4522 9454
rect 4556 9420 4590 9454
rect 4624 9420 4658 9454
rect 4692 9420 4726 9454
rect 4760 9420 4794 9454
rect 4828 9420 4862 9454
rect 4896 9420 4930 9454
rect 4964 9420 4998 9454
rect 5032 9420 5066 9454
rect 5100 9420 5134 9454
rect 5168 9420 5202 9454
rect 5236 9420 5270 9454
rect 5304 9420 5338 9454
rect 5372 9420 5406 9454
rect 5440 9420 5474 9454
rect 5508 9420 5542 9454
rect 5576 9420 5610 9454
rect 5644 9420 5678 9454
rect 5712 9420 5746 9454
rect 5780 9420 5814 9454
rect 5848 9420 5882 9454
rect 5916 9420 5950 9454
rect 5984 9420 6018 9454
rect 6052 9420 6086 9454
rect 6120 9420 6154 9454
rect 6188 9420 6222 9454
rect 6256 9420 6290 9454
rect 6324 9420 6358 9454
rect 6392 9420 6426 9454
rect 6460 9420 6494 9454
rect 6528 9420 6562 9454
rect 6596 9420 6630 9454
rect 6664 9420 6698 9454
rect 6732 9420 6766 9454
rect 6800 9420 6834 9454
rect 6868 9420 6902 9454
rect 6936 9420 6970 9454
rect 7004 9420 7038 9454
rect 7072 9420 7106 9454
rect 7140 9420 7174 9454
rect 7208 9420 7242 9454
rect 7276 9420 7310 9454
rect 7344 9420 7378 9454
rect 7412 9420 7446 9454
rect 7480 9420 7514 9454
rect 7548 9420 7582 9454
rect 7616 9420 7650 9454
rect 7684 9420 7718 9454
rect 7752 9420 7786 9454
rect 7820 9420 7854 9454
rect 7888 9420 7922 9454
rect 7956 9420 7990 9454
rect 8024 9420 8058 9454
rect 8092 9420 8126 9454
rect 8160 9420 8194 9454
rect 8228 9420 8262 9454
rect 8296 9420 8330 9454
rect 8364 9420 8398 9454
rect 8432 9420 8466 9454
rect 8500 9420 8534 9454
rect 8568 9420 8602 9454
rect 8636 9420 8670 9454
rect 8704 9420 8738 9454
rect 8772 9420 8806 9454
rect 8840 9420 8874 9454
rect 8908 9420 8942 9454
rect 8976 9420 9010 9454
rect 9044 9420 9078 9454
rect 9112 9420 9146 9454
rect 9180 9420 9214 9454
rect 9248 9420 9282 9454
rect 9316 9420 9350 9454
rect 9384 9420 9418 9454
rect 9452 9420 9486 9454
rect 9520 9420 9554 9454
rect 9588 9420 9622 9454
rect 9656 9420 9690 9454
rect 9724 9420 9758 9454
rect 9792 9420 9826 9454
rect 9860 9420 9894 9454
rect 9928 9420 9962 9454
rect 9996 9420 10030 9454
rect 10064 9420 10098 9454
rect 10132 9420 10166 9454
rect 10200 9420 10234 9454
rect 10268 9420 10302 9454
rect 10336 9420 10370 9454
rect 10404 9420 10438 9454
rect 10472 9420 10506 9454
rect 10540 9420 10574 9454
rect 10608 9420 10642 9454
rect 10676 9420 10710 9454
rect 10744 9420 10778 9454
rect 10812 9420 10846 9454
rect 10880 9420 10914 9454
rect 10948 9420 10982 9454
rect 11016 9420 11050 9454
rect 11084 9420 11118 9454
rect 11152 9420 11186 9454
rect 11220 9420 11254 9454
rect 11288 9420 11322 9454
rect 11356 9420 11390 9454
rect 11424 9420 11458 9454
rect 11492 9420 11526 9454
rect 11560 9420 11594 9454
rect 11628 9420 11662 9454
rect 11696 9420 11730 9454
rect 11764 9420 11798 9454
rect 11832 9420 11866 9454
rect 11900 9420 11934 9454
rect 11968 9420 12002 9454
rect 12036 9420 12070 9454
rect 12104 9420 12138 9454
rect 12172 9420 12206 9454
rect 12240 9420 12274 9454
rect 12308 9420 12342 9454
rect 12376 9420 12410 9454
rect 12444 9420 12478 9454
rect 12512 9420 12546 9454
rect 12580 9420 12614 9454
rect 12648 9420 12682 9454
rect 12716 9420 12750 9454
rect 12784 9420 12818 9454
rect 12852 9420 12886 9454
rect 12920 9420 12954 9454
rect 12988 9420 13022 9454
rect 13056 9420 13090 9454
rect 13124 9420 13158 9454
rect 13192 9420 13226 9454
rect 13260 9420 13294 9454
rect 13328 9420 13362 9454
rect 13396 9420 13430 9454
rect 13464 9420 13498 9454
rect 13532 9420 13566 9454
rect 13600 9420 13634 9454
rect 13668 9420 13702 9454
rect 13736 9420 13770 9454
rect 13804 9420 13838 9454
rect 13872 9420 13906 9454
rect 13940 9420 13974 9454
rect 14008 9420 14042 9454
rect 14076 9420 14110 9454
rect 14144 9420 14178 9454
rect 14212 9420 14246 9454
rect 14280 9420 14314 9454
rect 14348 9420 14382 9454
rect 14416 9420 14450 9454
rect 14484 9420 14724 9454
rect 245 9343 14724 9420
<< mvnsubdiff >>
rect 597 36177 14381 36227
rect 597 36143 773 36177
rect 807 36143 841 36177
rect 875 36143 909 36177
rect 943 36143 977 36177
rect 1011 36143 1045 36177
rect 1079 36143 1113 36177
rect 1147 36143 1181 36177
rect 1215 36143 1249 36177
rect 1283 36143 1317 36177
rect 1351 36143 1385 36177
rect 1419 36143 1453 36177
rect 1487 36143 1521 36177
rect 1555 36143 1589 36177
rect 1623 36143 1657 36177
rect 1691 36143 1725 36177
rect 1759 36143 1793 36177
rect 1827 36143 1861 36177
rect 1895 36143 1929 36177
rect 1963 36143 1997 36177
rect 2031 36143 2065 36177
rect 2099 36143 2133 36177
rect 2167 36143 2201 36177
rect 2235 36143 2269 36177
rect 2303 36143 2337 36177
rect 2371 36143 2405 36177
rect 2439 36143 2473 36177
rect 2507 36143 2541 36177
rect 2575 36143 2609 36177
rect 2643 36143 2677 36177
rect 2711 36143 2745 36177
rect 2779 36143 2813 36177
rect 2847 36143 2881 36177
rect 2915 36143 2949 36177
rect 2983 36143 3017 36177
rect 3051 36143 3085 36177
rect 3119 36143 3153 36177
rect 3187 36143 3221 36177
rect 3255 36143 3289 36177
rect 3323 36143 3357 36177
rect 3391 36143 3425 36177
rect 3459 36143 3493 36177
rect 3527 36143 3561 36177
rect 3595 36143 3629 36177
rect 3663 36143 3697 36177
rect 3731 36143 3765 36177
rect 3799 36143 3833 36177
rect 3867 36143 3901 36177
rect 3935 36143 3969 36177
rect 4003 36143 4037 36177
rect 4071 36143 4105 36177
rect 4139 36143 4173 36177
rect 4207 36143 4241 36177
rect 4275 36143 4309 36177
rect 4343 36143 4377 36177
rect 4411 36143 4445 36177
rect 4479 36143 4513 36177
rect 4547 36143 4581 36177
rect 4615 36143 4649 36177
rect 4683 36143 4717 36177
rect 4751 36143 4785 36177
rect 4819 36143 4853 36177
rect 4887 36143 4921 36177
rect 4955 36143 4989 36177
rect 5023 36143 5057 36177
rect 5091 36143 5125 36177
rect 5159 36143 5193 36177
rect 5227 36143 5261 36177
rect 5295 36143 5329 36177
rect 5363 36143 5397 36177
rect 5431 36143 5465 36177
rect 5499 36143 5533 36177
rect 5567 36143 5601 36177
rect 5635 36143 5669 36177
rect 5703 36143 5737 36177
rect 5771 36143 5805 36177
rect 5839 36143 5873 36177
rect 5907 36143 5941 36177
rect 5975 36143 6009 36177
rect 6043 36143 6077 36177
rect 6111 36143 6145 36177
rect 6179 36143 6213 36177
rect 6247 36143 6281 36177
rect 6315 36143 6349 36177
rect 6383 36143 6417 36177
rect 6451 36143 6485 36177
rect 6519 36143 6553 36177
rect 6587 36143 6621 36177
rect 6655 36143 6689 36177
rect 6723 36143 6757 36177
rect 6791 36143 6825 36177
rect 6859 36143 6893 36177
rect 6927 36143 6961 36177
rect 6995 36143 7029 36177
rect 7063 36143 7097 36177
rect 7131 36143 7165 36177
rect 7199 36143 7233 36177
rect 7267 36143 7301 36177
rect 7335 36143 7369 36177
rect 7403 36143 7437 36177
rect 7471 36143 7505 36177
rect 7539 36143 7573 36177
rect 7607 36143 7641 36177
rect 7675 36143 7709 36177
rect 7743 36143 7777 36177
rect 7811 36143 7845 36177
rect 7879 36143 7913 36177
rect 7947 36143 7981 36177
rect 8015 36143 8049 36177
rect 8083 36143 8117 36177
rect 8151 36143 8185 36177
rect 8219 36143 8253 36177
rect 8287 36143 8321 36177
rect 8355 36143 8389 36177
rect 8423 36143 8457 36177
rect 8491 36143 8525 36177
rect 8559 36143 8593 36177
rect 8627 36143 8661 36177
rect 8695 36143 8729 36177
rect 8763 36143 8797 36177
rect 8831 36143 8865 36177
rect 8899 36143 8933 36177
rect 8967 36143 9001 36177
rect 9035 36143 9069 36177
rect 9103 36143 9137 36177
rect 9171 36143 9205 36177
rect 9239 36143 9273 36177
rect 9307 36143 9341 36177
rect 9375 36143 9409 36177
rect 9443 36143 9477 36177
rect 9511 36143 9545 36177
rect 9579 36143 9613 36177
rect 9647 36143 9681 36177
rect 9715 36143 9749 36177
rect 9783 36143 9817 36177
rect 9851 36143 9885 36177
rect 9919 36143 9953 36177
rect 9987 36143 10021 36177
rect 10055 36143 10089 36177
rect 10123 36143 10157 36177
rect 10191 36143 10225 36177
rect 10259 36143 10293 36177
rect 10327 36143 10361 36177
rect 10395 36143 10429 36177
rect 10463 36143 10497 36177
rect 10531 36143 10565 36177
rect 10599 36143 10633 36177
rect 10667 36143 10701 36177
rect 10735 36143 10769 36177
rect 10803 36143 10837 36177
rect 10871 36143 10905 36177
rect 10939 36143 10973 36177
rect 11007 36143 11041 36177
rect 11075 36143 11109 36177
rect 11143 36143 11177 36177
rect 11211 36143 11245 36177
rect 11279 36143 11313 36177
rect 11347 36143 11381 36177
rect 11415 36143 11449 36177
rect 11483 36143 11517 36177
rect 11551 36143 11585 36177
rect 11619 36143 11653 36177
rect 11687 36143 11721 36177
rect 11755 36143 11789 36177
rect 11823 36143 11857 36177
rect 11891 36143 11925 36177
rect 11959 36143 11993 36177
rect 12027 36143 12061 36177
rect 12095 36143 12129 36177
rect 12163 36143 12197 36177
rect 12231 36143 12265 36177
rect 12299 36143 12333 36177
rect 12367 36143 12401 36177
rect 12435 36143 12469 36177
rect 12503 36143 12537 36177
rect 12571 36143 12605 36177
rect 12639 36143 12673 36177
rect 12707 36143 12741 36177
rect 12775 36143 12809 36177
rect 12843 36143 12877 36177
rect 12911 36143 12945 36177
rect 12979 36143 13013 36177
rect 13047 36143 13081 36177
rect 13115 36143 13149 36177
rect 13183 36143 13217 36177
rect 13251 36143 13285 36177
rect 13319 36143 13353 36177
rect 13387 36143 13421 36177
rect 13455 36143 13489 36177
rect 13523 36143 13557 36177
rect 13591 36143 13625 36177
rect 13659 36143 13693 36177
rect 13727 36143 13761 36177
rect 13795 36143 13829 36177
rect 13863 36143 13897 36177
rect 13931 36143 13965 36177
rect 13999 36143 14033 36177
rect 14067 36143 14101 36177
rect 14135 36143 14169 36177
rect 14203 36143 14381 36177
rect 597 36093 14381 36143
rect 597 36032 729 36093
rect 597 35998 646 36032
rect 680 35998 729 36032
rect 597 35964 729 35998
rect 597 35930 646 35964
rect 680 35930 729 35964
rect 597 35896 729 35930
rect 597 35862 646 35896
rect 680 35862 729 35896
rect 597 35828 729 35862
rect 597 35794 646 35828
rect 680 35794 729 35828
rect 597 35760 729 35794
rect 597 35726 646 35760
rect 680 35726 729 35760
rect 597 35692 729 35726
rect 597 35658 646 35692
rect 680 35658 729 35692
rect 597 35624 729 35658
rect 597 35590 646 35624
rect 680 35590 729 35624
rect 597 35556 729 35590
rect 597 35522 646 35556
rect 680 35522 729 35556
rect 597 35488 729 35522
rect 597 35454 646 35488
rect 680 35454 729 35488
rect 597 35420 729 35454
rect 597 35386 646 35420
rect 680 35386 729 35420
rect 597 35352 729 35386
rect 597 35318 646 35352
rect 680 35318 729 35352
rect 597 35284 729 35318
rect 597 35250 646 35284
rect 680 35250 729 35284
rect 597 35216 729 35250
rect 597 35182 646 35216
rect 680 35182 729 35216
rect 597 35148 729 35182
rect 597 35114 646 35148
rect 680 35114 729 35148
rect 597 35080 729 35114
rect 597 35046 646 35080
rect 680 35046 729 35080
rect 597 35012 729 35046
rect 597 34978 646 35012
rect 680 34978 729 35012
rect 597 34944 729 34978
rect 597 34910 646 34944
rect 680 34910 729 34944
rect 597 34876 729 34910
rect 597 34842 646 34876
rect 680 34842 729 34876
rect 597 34808 729 34842
rect 597 34774 646 34808
rect 680 34774 729 34808
rect 597 34740 729 34774
rect 597 34706 646 34740
rect 680 34706 729 34740
rect 597 34672 729 34706
rect 14247 36032 14381 36093
rect 14247 35998 14297 36032
rect 14331 35998 14381 36032
rect 14247 35964 14381 35998
rect 14247 35930 14297 35964
rect 14331 35930 14381 35964
rect 14247 35896 14381 35930
rect 14247 35862 14297 35896
rect 14331 35862 14381 35896
rect 14247 35828 14381 35862
rect 14247 35794 14297 35828
rect 14331 35794 14381 35828
rect 14247 35760 14381 35794
rect 14247 35726 14297 35760
rect 14331 35726 14381 35760
rect 14247 35692 14381 35726
rect 14247 35658 14297 35692
rect 14331 35658 14381 35692
rect 14247 35624 14381 35658
rect 14247 35590 14297 35624
rect 14331 35590 14381 35624
rect 14247 35556 14381 35590
rect 14247 35522 14297 35556
rect 14331 35522 14381 35556
rect 14247 35488 14381 35522
rect 14247 35454 14297 35488
rect 14331 35454 14381 35488
rect 14247 35420 14381 35454
rect 14247 35386 14297 35420
rect 14331 35386 14381 35420
rect 14247 35352 14381 35386
rect 14247 35318 14297 35352
rect 14331 35318 14381 35352
rect 14247 35284 14381 35318
rect 14247 35250 14297 35284
rect 14331 35250 14381 35284
rect 14247 35216 14381 35250
rect 14247 35182 14297 35216
rect 14331 35182 14381 35216
rect 14247 35148 14381 35182
rect 14247 35114 14297 35148
rect 14331 35114 14381 35148
rect 14247 35080 14381 35114
rect 14247 35046 14297 35080
rect 14331 35046 14381 35080
rect 14247 35012 14381 35046
rect 14247 34978 14297 35012
rect 14331 34978 14381 35012
rect 14247 34944 14381 34978
rect 14247 34910 14297 34944
rect 14331 34910 14381 34944
rect 14247 34876 14381 34910
rect 14247 34842 14297 34876
rect 14331 34842 14381 34876
rect 14247 34808 14381 34842
rect 14247 34774 14297 34808
rect 14331 34774 14381 34808
rect 14247 34740 14381 34774
rect 14247 34706 14297 34740
rect 14331 34706 14381 34740
rect 597 34638 646 34672
rect 680 34638 729 34672
rect 597 34604 729 34638
rect 597 34570 646 34604
rect 680 34570 729 34604
rect 597 34536 729 34570
rect 597 34502 646 34536
rect 680 34502 729 34536
rect 597 34468 729 34502
rect 597 34434 646 34468
rect 680 34434 729 34468
rect 597 34400 729 34434
rect 597 34366 646 34400
rect 680 34366 729 34400
rect 597 34332 729 34366
rect 597 34298 646 34332
rect 680 34298 729 34332
rect 597 34264 729 34298
rect 597 34230 646 34264
rect 680 34230 729 34264
rect 597 34196 729 34230
rect 597 34162 646 34196
rect 680 34162 729 34196
rect 597 34128 729 34162
rect 597 34094 646 34128
rect 680 34094 729 34128
rect 597 34060 729 34094
rect 597 34026 646 34060
rect 680 34026 729 34060
rect 597 33992 729 34026
rect 597 33958 646 33992
rect 680 33958 729 33992
rect 597 33924 729 33958
rect 597 33890 646 33924
rect 680 33890 729 33924
rect 597 33856 729 33890
rect 597 33822 646 33856
rect 680 33822 729 33856
rect 597 33788 729 33822
rect 597 33754 646 33788
rect 680 33754 729 33788
rect 597 33720 729 33754
rect 597 33686 646 33720
rect 680 33686 729 33720
rect 597 33652 729 33686
rect 597 33618 646 33652
rect 680 33618 729 33652
rect 597 33584 729 33618
rect 597 33550 646 33584
rect 680 33550 729 33584
rect 597 33516 729 33550
rect 597 33482 646 33516
rect 680 33482 729 33516
rect 597 33448 729 33482
rect 597 33414 646 33448
rect 680 33414 729 33448
rect 597 33380 729 33414
rect 597 33346 646 33380
rect 680 33346 729 33380
rect 597 33312 729 33346
rect 597 33278 646 33312
rect 680 33278 729 33312
rect 597 33244 729 33278
rect 597 33210 646 33244
rect 680 33210 729 33244
rect 597 33176 729 33210
rect 597 33142 646 33176
rect 680 33142 729 33176
rect 597 33108 729 33142
rect 597 33074 646 33108
rect 680 33074 729 33108
rect 597 33040 729 33074
rect 597 33006 646 33040
rect 680 33006 729 33040
rect 597 32972 729 33006
rect 597 32938 646 32972
rect 680 32938 729 32972
rect 597 32904 729 32938
rect 597 32870 646 32904
rect 680 32870 729 32904
rect 597 32836 729 32870
rect 597 32802 646 32836
rect 680 32802 729 32836
rect 597 32768 729 32802
rect 597 32734 646 32768
rect 680 32734 729 32768
rect 597 32700 729 32734
rect 597 32666 646 32700
rect 680 32666 729 32700
rect 597 32632 729 32666
rect 597 32598 646 32632
rect 680 32598 729 32632
rect 597 32564 729 32598
rect 597 32530 646 32564
rect 680 32530 729 32564
rect 597 32496 729 32530
rect 597 32462 646 32496
rect 680 32462 729 32496
rect 597 32428 729 32462
rect 597 32394 646 32428
rect 680 32394 729 32428
rect 597 32360 729 32394
rect 597 32326 646 32360
rect 680 32326 729 32360
rect 597 32292 729 32326
rect 597 32258 646 32292
rect 680 32258 729 32292
rect 597 32224 729 32258
rect 597 32190 646 32224
rect 680 32190 729 32224
rect 597 32156 729 32190
rect 597 32122 646 32156
rect 680 32122 729 32156
rect 597 32088 729 32122
rect 597 32054 646 32088
rect 680 32054 729 32088
rect 597 32020 729 32054
rect 597 31986 646 32020
rect 680 31986 729 32020
rect 597 31952 729 31986
rect 597 31918 646 31952
rect 680 31918 729 31952
rect 597 31884 729 31918
rect 597 31850 646 31884
rect 680 31850 729 31884
rect 597 31816 729 31850
rect 597 31782 646 31816
rect 680 31782 729 31816
rect 597 31748 729 31782
rect 597 31714 646 31748
rect 680 31714 729 31748
rect 597 31680 729 31714
rect 597 31646 646 31680
rect 680 31646 729 31680
rect 597 31612 729 31646
rect 597 31578 646 31612
rect 680 31578 729 31612
rect 597 31544 729 31578
rect 597 31510 646 31544
rect 680 31510 729 31544
rect 597 31476 729 31510
rect 597 31442 646 31476
rect 680 31442 729 31476
rect 597 31408 729 31442
rect 597 31374 646 31408
rect 680 31374 729 31408
rect 597 31340 729 31374
rect 597 31306 646 31340
rect 680 31306 729 31340
rect 597 31272 729 31306
rect 597 31238 646 31272
rect 680 31238 729 31272
rect 597 31204 729 31238
rect 597 31170 646 31204
rect 680 31170 729 31204
rect 597 31136 729 31170
rect 597 31102 646 31136
rect 680 31102 729 31136
rect 597 31068 729 31102
rect 597 31034 646 31068
rect 680 31034 729 31068
rect 597 31000 729 31034
rect 597 30966 646 31000
rect 680 30966 729 31000
rect 597 30932 729 30966
rect 597 30898 646 30932
rect 680 30898 729 30932
rect 597 30864 729 30898
rect 597 30830 646 30864
rect 680 30830 729 30864
rect 597 30796 729 30830
rect 597 30762 646 30796
rect 680 30762 729 30796
rect 597 30728 729 30762
rect 597 30694 646 30728
rect 680 30694 729 30728
rect 597 30660 729 30694
rect 597 30626 646 30660
rect 680 30626 729 30660
rect 597 30592 729 30626
rect 597 30558 646 30592
rect 680 30558 729 30592
rect 597 30524 729 30558
rect 597 30490 646 30524
rect 680 30490 729 30524
rect 597 30456 729 30490
rect 597 30422 646 30456
rect 680 30422 729 30456
rect 597 30388 729 30422
rect 597 30354 646 30388
rect 680 30354 729 30388
rect 597 30320 729 30354
rect 597 30286 646 30320
rect 680 30286 729 30320
rect 597 30252 729 30286
rect 597 30218 646 30252
rect 680 30218 729 30252
rect 597 30184 729 30218
rect 597 30150 646 30184
rect 680 30150 729 30184
rect 597 30116 729 30150
rect 597 30082 646 30116
rect 680 30082 729 30116
rect 597 30048 729 30082
rect 597 30014 646 30048
rect 680 30014 729 30048
rect 597 29980 729 30014
rect 597 29946 646 29980
rect 680 29946 729 29980
rect 597 29912 729 29946
rect 597 29878 646 29912
rect 680 29878 729 29912
rect 597 29844 729 29878
rect 597 29810 646 29844
rect 680 29810 729 29844
rect 597 29776 729 29810
rect 597 29742 646 29776
rect 680 29742 729 29776
rect 597 29708 729 29742
rect 597 29674 646 29708
rect 680 29674 729 29708
rect 597 29640 729 29674
rect 597 29606 646 29640
rect 680 29606 729 29640
rect 597 29572 729 29606
rect 597 29538 646 29572
rect 680 29538 729 29572
rect 597 29504 729 29538
rect 597 29470 646 29504
rect 680 29470 729 29504
rect 597 29436 729 29470
rect 597 29402 646 29436
rect 680 29402 729 29436
rect 597 29368 729 29402
rect 597 29334 646 29368
rect 680 29334 729 29368
rect 597 29300 729 29334
rect 597 29266 646 29300
rect 680 29266 729 29300
rect 597 29232 729 29266
rect 597 29198 646 29232
rect 680 29198 729 29232
rect 597 29164 729 29198
rect 597 29130 646 29164
rect 680 29130 729 29164
rect 597 29096 729 29130
rect 597 29062 646 29096
rect 680 29062 729 29096
rect 597 29028 729 29062
rect 597 28994 646 29028
rect 680 28994 729 29028
rect 597 28960 729 28994
rect 597 28926 646 28960
rect 680 28926 729 28960
rect 597 28892 729 28926
rect 597 28858 646 28892
rect 680 28858 729 28892
rect 597 28824 729 28858
rect 597 28790 646 28824
rect 680 28790 729 28824
rect 597 28756 729 28790
rect 597 28722 646 28756
rect 680 28722 729 28756
rect 597 28688 729 28722
rect 597 28654 646 28688
rect 680 28654 729 28688
rect 597 28620 729 28654
rect 597 28586 646 28620
rect 680 28586 729 28620
rect 597 28552 729 28586
rect 597 28518 646 28552
rect 680 28518 729 28552
rect 597 28484 729 28518
rect 597 28450 646 28484
rect 680 28450 729 28484
rect 597 28416 729 28450
rect 597 28382 646 28416
rect 680 28382 729 28416
rect 597 28348 729 28382
rect 597 28314 646 28348
rect 680 28314 729 28348
rect 597 28280 729 28314
rect 597 28246 646 28280
rect 680 28246 729 28280
rect 597 28212 729 28246
rect 597 28178 646 28212
rect 680 28178 729 28212
rect 597 28144 729 28178
rect 597 28110 646 28144
rect 680 28110 729 28144
rect 597 28076 729 28110
rect 597 28042 646 28076
rect 680 28042 729 28076
rect 597 28008 729 28042
rect 597 27974 646 28008
rect 680 27974 729 28008
rect 597 27940 729 27974
rect 597 27906 646 27940
rect 680 27906 729 27940
rect 597 27872 729 27906
rect 597 27838 646 27872
rect 680 27838 729 27872
rect 597 27804 729 27838
rect 597 27770 646 27804
rect 680 27770 729 27804
rect 597 27736 729 27770
rect 597 27702 646 27736
rect 680 27702 729 27736
rect 597 27668 729 27702
rect 597 27634 646 27668
rect 680 27634 729 27668
rect 597 27600 729 27634
rect 597 27566 646 27600
rect 680 27566 729 27600
rect 597 27532 729 27566
rect 597 27498 646 27532
rect 680 27498 729 27532
rect 597 27464 729 27498
rect 597 27430 646 27464
rect 680 27430 729 27464
rect 597 27396 729 27430
rect 597 27362 646 27396
rect 680 27362 729 27396
rect 597 27328 729 27362
rect 597 27294 646 27328
rect 680 27294 729 27328
rect 597 27260 729 27294
rect 597 27226 646 27260
rect 680 27226 729 27260
rect 597 27192 729 27226
rect 597 27158 646 27192
rect 680 27158 729 27192
rect 597 27124 729 27158
rect 597 27090 646 27124
rect 680 27090 729 27124
rect 597 27056 729 27090
rect 597 27022 646 27056
rect 680 27022 729 27056
rect 597 26988 729 27022
rect 597 26954 646 26988
rect 680 26954 729 26988
rect 597 26920 729 26954
rect 597 26886 646 26920
rect 680 26886 729 26920
rect 597 26852 729 26886
rect 597 26818 646 26852
rect 680 26818 729 26852
rect 597 26784 729 26818
rect 597 26750 646 26784
rect 680 26750 729 26784
rect 597 26716 729 26750
rect 597 26682 646 26716
rect 680 26682 729 26716
rect 597 26648 729 26682
rect 597 26614 646 26648
rect 680 26614 729 26648
rect 597 26580 729 26614
rect 597 26546 646 26580
rect 680 26546 729 26580
rect 597 26512 729 26546
rect 597 26478 646 26512
rect 680 26478 729 26512
rect 597 26444 729 26478
rect 597 26410 646 26444
rect 680 26410 729 26444
rect 597 26376 729 26410
rect 597 26342 646 26376
rect 680 26342 729 26376
rect 597 26308 729 26342
rect 597 26274 646 26308
rect 680 26274 729 26308
rect 597 26240 729 26274
rect 597 26206 646 26240
rect 680 26206 729 26240
rect 597 26172 729 26206
rect 597 26138 646 26172
rect 680 26138 729 26172
rect 597 26104 729 26138
rect 597 26070 646 26104
rect 680 26070 729 26104
rect 597 26036 729 26070
rect 597 26002 646 26036
rect 680 26002 729 26036
rect 597 25968 729 26002
rect 597 25934 646 25968
rect 680 25934 729 25968
rect 597 25900 729 25934
rect 597 25866 646 25900
rect 680 25866 729 25900
rect 597 25832 729 25866
rect 597 25798 646 25832
rect 680 25798 729 25832
rect 597 25764 729 25798
rect 597 25730 646 25764
rect 680 25730 729 25764
rect 597 25696 729 25730
rect 597 25662 646 25696
rect 680 25662 729 25696
rect 597 25628 729 25662
rect 597 25594 646 25628
rect 680 25594 729 25628
rect 597 25560 729 25594
rect 597 25526 646 25560
rect 680 25526 729 25560
rect 597 25492 729 25526
rect 597 25458 646 25492
rect 680 25458 729 25492
rect 597 25424 729 25458
rect 597 25390 646 25424
rect 680 25390 729 25424
rect 597 25356 729 25390
rect 597 25322 646 25356
rect 680 25322 729 25356
rect 597 25288 729 25322
rect 597 25254 646 25288
rect 680 25254 729 25288
rect 597 25220 729 25254
rect 597 25186 646 25220
rect 680 25186 729 25220
rect 597 25152 729 25186
rect 597 25118 646 25152
rect 680 25118 729 25152
rect 597 25084 729 25118
rect 597 25050 646 25084
rect 680 25050 729 25084
rect 597 25016 729 25050
rect 597 24982 646 25016
rect 680 24982 729 25016
rect 597 24948 729 24982
rect 597 24914 646 24948
rect 680 24914 729 24948
rect 597 24880 729 24914
rect 597 24846 646 24880
rect 680 24846 729 24880
rect 597 24812 729 24846
rect 597 24778 646 24812
rect 680 24778 729 24812
rect 597 24744 729 24778
rect 597 24710 646 24744
rect 680 24710 729 24744
rect 597 24676 729 24710
rect 597 24642 646 24676
rect 680 24642 729 24676
rect 597 24608 729 24642
rect 597 24574 646 24608
rect 680 24574 729 24608
rect 597 24540 729 24574
rect 597 24506 646 24540
rect 680 24506 729 24540
rect 597 24472 729 24506
rect 597 24438 646 24472
rect 680 24438 729 24472
rect 597 24404 729 24438
rect 597 24370 646 24404
rect 680 24370 729 24404
rect 597 24336 729 24370
rect 597 24302 646 24336
rect 680 24302 729 24336
rect 597 24268 729 24302
rect 597 24234 646 24268
rect 680 24234 729 24268
rect 597 24200 729 24234
rect 597 24166 646 24200
rect 680 24166 729 24200
rect 597 24132 729 24166
rect 597 24098 646 24132
rect 680 24098 729 24132
rect 597 24064 729 24098
rect 597 24030 646 24064
rect 680 24030 729 24064
rect 597 23996 729 24030
rect 597 23962 646 23996
rect 680 23962 729 23996
rect 597 23928 729 23962
rect 597 23894 646 23928
rect 680 23894 729 23928
rect 597 23860 729 23894
rect 597 23826 646 23860
rect 680 23826 729 23860
rect 597 23792 729 23826
rect 597 23758 646 23792
rect 680 23758 729 23792
rect 597 23724 729 23758
rect 597 23690 646 23724
rect 680 23690 729 23724
rect 597 23656 729 23690
rect 597 23622 646 23656
rect 680 23622 729 23656
rect 597 23588 729 23622
rect 597 23554 646 23588
rect 680 23554 729 23588
rect 597 23520 729 23554
rect 597 23486 646 23520
rect 680 23486 729 23520
rect 597 23452 729 23486
rect 597 23418 646 23452
rect 680 23418 729 23452
rect 597 23384 729 23418
rect 597 23350 646 23384
rect 680 23350 729 23384
rect 597 23316 729 23350
rect 597 23282 646 23316
rect 680 23282 729 23316
rect 597 23248 729 23282
rect 597 23214 646 23248
rect 680 23214 729 23248
rect 597 23180 729 23214
rect 597 23146 646 23180
rect 680 23146 729 23180
rect 597 23112 729 23146
rect 597 23078 646 23112
rect 680 23078 729 23112
rect 597 23044 729 23078
rect 597 23010 646 23044
rect 680 23010 729 23044
rect 597 22976 729 23010
rect 597 22942 646 22976
rect 680 22942 729 22976
rect 597 22908 729 22942
rect 597 22874 646 22908
rect 680 22874 729 22908
rect 597 22840 729 22874
rect 597 22806 646 22840
rect 680 22806 729 22840
rect 597 22772 729 22806
rect 597 22738 646 22772
rect 680 22738 729 22772
rect 597 22704 729 22738
rect 597 22670 646 22704
rect 680 22670 729 22704
rect 597 22636 729 22670
rect 597 22602 646 22636
rect 680 22602 729 22636
rect 597 22568 729 22602
rect 597 22534 646 22568
rect 680 22534 729 22568
rect 597 22500 729 22534
rect 597 22466 646 22500
rect 680 22466 729 22500
rect 597 22432 729 22466
rect 597 22398 646 22432
rect 680 22398 729 22432
rect 597 22364 729 22398
rect 597 22330 646 22364
rect 680 22330 729 22364
rect 597 22296 729 22330
rect 597 22262 646 22296
rect 680 22262 729 22296
rect 597 22228 729 22262
rect 597 22194 646 22228
rect 680 22194 729 22228
rect 597 22160 729 22194
rect 597 22126 646 22160
rect 680 22126 729 22160
rect 597 22092 729 22126
rect 597 22058 646 22092
rect 680 22058 729 22092
rect 597 22024 729 22058
rect 597 21990 646 22024
rect 680 21990 729 22024
rect 597 21956 729 21990
rect 597 21922 646 21956
rect 680 21922 729 21956
rect 597 21888 729 21922
rect 597 21854 646 21888
rect 680 21854 729 21888
rect 597 21820 729 21854
rect 597 21786 646 21820
rect 680 21786 729 21820
rect 597 21752 729 21786
rect 597 21718 646 21752
rect 680 21718 729 21752
rect 597 21684 729 21718
rect 597 21650 646 21684
rect 680 21650 729 21684
rect 597 21616 729 21650
rect 597 21582 646 21616
rect 680 21582 729 21616
rect 597 21548 729 21582
rect 597 21514 646 21548
rect 680 21514 729 21548
rect 597 21480 729 21514
rect 597 21446 646 21480
rect 680 21446 729 21480
rect 597 21412 729 21446
rect 597 21378 646 21412
rect 680 21378 729 21412
rect 597 21344 729 21378
rect 597 21310 646 21344
rect 680 21310 729 21344
rect 597 21276 729 21310
rect 597 21242 646 21276
rect 680 21242 729 21276
rect 597 21208 729 21242
rect 597 21174 646 21208
rect 680 21174 729 21208
rect 597 21140 729 21174
rect 597 21106 646 21140
rect 680 21106 729 21140
rect 597 21072 729 21106
rect 597 21038 646 21072
rect 680 21038 729 21072
rect 597 21004 729 21038
rect 597 20970 646 21004
rect 680 20970 729 21004
rect 597 20936 729 20970
rect 597 20902 646 20936
rect 680 20902 729 20936
rect 597 20868 729 20902
rect 597 20834 646 20868
rect 680 20834 729 20868
rect 597 20800 729 20834
rect 597 20766 646 20800
rect 680 20766 729 20800
rect 597 20732 729 20766
rect 597 20698 646 20732
rect 680 20698 729 20732
rect 597 20664 729 20698
rect 597 20630 646 20664
rect 680 20630 729 20664
rect 597 20596 729 20630
rect 597 20562 646 20596
rect 680 20562 729 20596
rect 597 20528 729 20562
rect 597 20494 646 20528
rect 680 20494 729 20528
rect 597 20460 729 20494
rect 597 20426 646 20460
rect 680 20426 729 20460
rect 597 20392 729 20426
rect 597 20358 646 20392
rect 680 20358 729 20392
rect 597 20324 729 20358
rect 597 20290 646 20324
rect 680 20290 729 20324
rect 597 20256 729 20290
rect 597 20222 646 20256
rect 680 20222 729 20256
rect 597 20188 729 20222
rect 597 20154 646 20188
rect 680 20154 729 20188
rect 597 20120 729 20154
rect 597 20086 646 20120
rect 680 20086 729 20120
rect 597 20052 729 20086
rect 597 20018 646 20052
rect 680 20018 729 20052
rect 597 19984 729 20018
rect 597 19950 646 19984
rect 680 19950 729 19984
rect 597 19916 729 19950
rect 597 19882 646 19916
rect 680 19882 729 19916
rect 597 19848 729 19882
rect 597 19814 646 19848
rect 680 19814 729 19848
rect 597 19780 729 19814
rect 597 19746 646 19780
rect 680 19746 729 19780
rect 597 19712 729 19746
rect 597 19678 646 19712
rect 680 19678 729 19712
rect 597 19644 729 19678
rect 597 19610 646 19644
rect 680 19610 729 19644
rect 597 19576 729 19610
rect 597 19542 646 19576
rect 680 19542 729 19576
rect 597 19508 729 19542
rect 597 19474 646 19508
rect 680 19474 729 19508
rect 597 19440 729 19474
rect 597 19406 646 19440
rect 680 19406 729 19440
rect 597 19372 729 19406
rect 597 19338 646 19372
rect 680 19338 729 19372
rect 597 19304 729 19338
rect 597 19270 646 19304
rect 680 19270 729 19304
rect 597 19236 729 19270
rect 597 19202 646 19236
rect 680 19202 729 19236
rect 597 19168 729 19202
rect 597 19134 646 19168
rect 680 19134 729 19168
rect 597 19100 729 19134
rect 597 19066 646 19100
rect 680 19066 729 19100
rect 597 19032 729 19066
rect 597 18998 646 19032
rect 680 18998 729 19032
rect 597 18964 729 18998
rect 597 18930 646 18964
rect 680 18930 729 18964
rect 597 18896 729 18930
rect 597 18862 646 18896
rect 680 18862 729 18896
rect 597 18828 729 18862
rect 597 18794 646 18828
rect 680 18794 729 18828
rect 597 18760 729 18794
rect 597 18726 646 18760
rect 680 18726 729 18760
rect 597 18692 729 18726
rect 597 18658 646 18692
rect 680 18658 729 18692
rect 597 18624 729 18658
rect 597 18590 646 18624
rect 680 18590 729 18624
rect 597 18556 729 18590
rect 597 18522 646 18556
rect 680 18522 729 18556
rect 597 18488 729 18522
rect 597 18454 646 18488
rect 680 18454 729 18488
rect 597 18420 729 18454
rect 597 18386 646 18420
rect 680 18386 729 18420
rect 597 18352 729 18386
rect 597 18318 646 18352
rect 680 18318 729 18352
rect 597 18284 729 18318
rect 597 18250 646 18284
rect 680 18250 729 18284
rect 597 18216 729 18250
rect 597 18182 646 18216
rect 680 18182 729 18216
rect 597 18148 729 18182
rect 597 18114 646 18148
rect 680 18114 729 18148
rect 597 18080 729 18114
rect 597 18046 646 18080
rect 680 18046 729 18080
rect 597 18012 729 18046
rect 597 17978 646 18012
rect 680 17978 729 18012
rect 597 17944 729 17978
rect 597 17910 646 17944
rect 680 17910 729 17944
rect 597 17876 729 17910
rect 597 17842 646 17876
rect 680 17842 729 17876
rect 597 17808 729 17842
rect 597 17774 646 17808
rect 680 17774 729 17808
rect 597 17740 729 17774
rect 597 17706 646 17740
rect 680 17706 729 17740
rect 597 17672 729 17706
rect 597 17638 646 17672
rect 680 17638 729 17672
rect 597 17604 729 17638
rect 597 17570 646 17604
rect 680 17570 729 17604
rect 597 17536 729 17570
rect 597 17502 646 17536
rect 680 17502 729 17536
rect 597 17468 729 17502
rect 597 17434 646 17468
rect 680 17434 729 17468
rect 597 17400 729 17434
rect 597 17366 646 17400
rect 680 17366 729 17400
rect 597 17332 729 17366
rect 597 17298 646 17332
rect 680 17298 729 17332
rect 597 17264 729 17298
rect 597 17230 646 17264
rect 680 17230 729 17264
rect 597 17196 729 17230
rect 597 17162 646 17196
rect 680 17162 729 17196
rect 597 17128 729 17162
rect 597 17094 646 17128
rect 680 17094 729 17128
rect 597 17060 729 17094
rect 597 17026 646 17060
rect 680 17026 729 17060
rect 597 16992 729 17026
rect 597 16958 646 16992
rect 680 16958 729 16992
rect 597 16924 729 16958
rect 597 16890 646 16924
rect 680 16890 729 16924
rect 597 16856 729 16890
rect 597 16822 646 16856
rect 680 16822 729 16856
rect 597 16788 729 16822
rect 597 16754 646 16788
rect 680 16754 729 16788
rect 597 16720 729 16754
rect 597 16686 646 16720
rect 680 16686 729 16720
rect 597 16652 729 16686
rect 597 16618 646 16652
rect 680 16618 729 16652
rect 597 16584 729 16618
rect 597 16550 646 16584
rect 680 16550 729 16584
rect 597 16516 729 16550
rect 597 16482 646 16516
rect 680 16482 729 16516
rect 597 16448 729 16482
rect 597 16414 646 16448
rect 680 16414 729 16448
rect 597 16380 729 16414
rect 597 16346 646 16380
rect 680 16346 729 16380
rect 597 16312 729 16346
rect 597 16278 646 16312
rect 680 16278 729 16312
rect 597 16244 729 16278
rect 597 16210 646 16244
rect 680 16210 729 16244
rect 597 16176 729 16210
rect 597 16142 646 16176
rect 680 16142 729 16176
rect 597 16108 729 16142
rect 597 16074 646 16108
rect 680 16074 729 16108
rect 597 16040 729 16074
rect 597 16006 646 16040
rect 680 16006 729 16040
rect 597 15972 729 16006
rect 597 15938 646 15972
rect 680 15938 729 15972
rect 597 15904 729 15938
rect 597 15870 646 15904
rect 680 15870 729 15904
rect 597 15836 729 15870
rect 597 15802 646 15836
rect 680 15802 729 15836
rect 597 15768 729 15802
rect 597 15734 646 15768
rect 680 15734 729 15768
rect 597 15700 729 15734
rect 597 15666 646 15700
rect 680 15666 729 15700
rect 597 15632 729 15666
rect 597 15598 646 15632
rect 680 15598 729 15632
rect 597 15564 729 15598
rect 597 15530 646 15564
rect 680 15530 729 15564
rect 597 15496 729 15530
rect 597 15462 646 15496
rect 680 15462 729 15496
rect 597 15428 729 15462
rect 597 15394 646 15428
rect 680 15394 729 15428
rect 597 15360 729 15394
rect 597 15326 646 15360
rect 680 15326 729 15360
rect 597 15292 729 15326
rect 597 15258 646 15292
rect 680 15258 729 15292
rect 597 15224 729 15258
rect 597 15190 646 15224
rect 680 15190 729 15224
rect 597 15156 729 15190
rect 597 15122 646 15156
rect 680 15122 729 15156
rect 597 15088 729 15122
rect 597 15054 646 15088
rect 680 15054 729 15088
rect 597 15020 729 15054
rect 597 14986 646 15020
rect 680 14986 729 15020
rect 597 14952 729 14986
rect 597 14918 646 14952
rect 680 14918 729 14952
rect 597 14884 729 14918
rect 597 14850 646 14884
rect 680 14850 729 14884
rect 597 14816 729 14850
rect 597 14782 646 14816
rect 680 14782 729 14816
rect 597 14748 729 14782
rect 597 14714 646 14748
rect 680 14714 729 14748
rect 597 14680 729 14714
rect 597 14646 646 14680
rect 680 14646 729 14680
rect 597 14612 729 14646
rect 597 14578 646 14612
rect 680 14578 729 14612
rect 597 14544 729 14578
rect 597 14510 646 14544
rect 680 14510 729 14544
rect 597 14476 729 14510
rect 597 14442 646 14476
rect 680 14442 729 14476
rect 597 14408 729 14442
rect 597 14374 646 14408
rect 680 14374 729 14408
rect 597 14340 729 14374
rect 597 14306 646 14340
rect 680 14306 729 14340
rect 597 14272 729 14306
rect 597 14238 646 14272
rect 680 14238 729 14272
rect 597 14204 729 14238
rect 597 14170 646 14204
rect 680 14170 729 14204
rect 597 14136 729 14170
rect 597 14102 646 14136
rect 680 14102 729 14136
rect 597 14068 729 14102
rect 597 14034 646 14068
rect 680 14034 729 14068
rect 597 14000 729 14034
rect 597 13966 646 14000
rect 680 13966 729 14000
rect 597 13932 729 13966
rect 597 13898 646 13932
rect 680 13898 729 13932
rect 597 13864 729 13898
rect 597 13830 646 13864
rect 680 13830 729 13864
rect 597 13796 729 13830
rect 597 13762 646 13796
rect 680 13762 729 13796
rect 597 13728 729 13762
rect 597 13694 646 13728
rect 680 13694 729 13728
rect 597 13660 729 13694
rect 597 13626 646 13660
rect 680 13626 729 13660
rect 597 13592 729 13626
rect 597 13558 646 13592
rect 680 13558 729 13592
rect 597 13524 729 13558
rect 597 13490 646 13524
rect 680 13490 729 13524
rect 597 13456 729 13490
rect 597 13422 646 13456
rect 680 13422 729 13456
rect 597 13388 729 13422
rect 597 13354 646 13388
rect 680 13354 729 13388
rect 597 13320 729 13354
rect 597 13286 646 13320
rect 680 13286 729 13320
rect 597 13252 729 13286
rect 597 13218 646 13252
rect 680 13218 729 13252
rect 597 13184 729 13218
rect 597 13150 646 13184
rect 680 13150 729 13184
rect 597 13116 729 13150
rect 597 13082 646 13116
rect 680 13082 729 13116
rect 597 13048 729 13082
rect 597 13014 646 13048
rect 680 13014 729 13048
rect 597 12980 729 13014
rect 597 12946 646 12980
rect 680 12946 729 12980
rect 597 12912 729 12946
rect 597 12878 646 12912
rect 680 12878 729 12912
rect 597 12844 729 12878
rect 597 12810 646 12844
rect 680 12810 729 12844
rect 597 12776 729 12810
rect 597 12742 646 12776
rect 680 12742 729 12776
rect 597 12708 729 12742
rect 597 12674 646 12708
rect 680 12674 729 12708
rect 597 12640 729 12674
rect 597 12606 646 12640
rect 680 12606 729 12640
rect 597 12572 729 12606
rect 597 12538 646 12572
rect 680 12538 729 12572
rect 597 12504 729 12538
rect 597 12470 646 12504
rect 680 12470 729 12504
rect 597 12436 729 12470
rect 597 12402 646 12436
rect 680 12402 729 12436
rect 597 12368 729 12402
rect 597 12334 646 12368
rect 680 12334 729 12368
rect 597 12300 729 12334
rect 597 12266 646 12300
rect 680 12266 729 12300
rect 597 12232 729 12266
rect 597 12198 646 12232
rect 680 12198 729 12232
rect 597 12164 729 12198
rect 597 12130 646 12164
rect 680 12130 729 12164
rect 597 12096 729 12130
rect 597 12062 646 12096
rect 680 12062 729 12096
rect 597 12028 729 12062
rect 597 11994 646 12028
rect 680 11994 729 12028
rect 597 11960 729 11994
rect 597 11926 646 11960
rect 680 11926 729 11960
rect 597 11892 729 11926
rect 597 11858 646 11892
rect 680 11858 729 11892
rect 597 11824 729 11858
rect 597 11790 646 11824
rect 680 11790 729 11824
rect 597 11756 729 11790
rect 597 11722 646 11756
rect 680 11722 729 11756
rect 597 11688 729 11722
rect 597 11654 646 11688
rect 680 11654 729 11688
rect 597 11620 729 11654
rect 597 11586 646 11620
rect 680 11586 729 11620
rect 597 11552 729 11586
rect 597 11518 646 11552
rect 680 11518 729 11552
rect 597 11484 729 11518
rect 597 11450 646 11484
rect 680 11450 729 11484
rect 597 11416 729 11450
rect 597 11382 646 11416
rect 680 11382 729 11416
rect 597 11348 729 11382
rect 597 11314 646 11348
rect 680 11314 729 11348
rect 597 11280 729 11314
rect 597 11246 646 11280
rect 680 11246 729 11280
rect 597 11212 729 11246
rect 597 11178 646 11212
rect 680 11178 729 11212
rect 597 11144 729 11178
rect 597 11110 646 11144
rect 680 11110 729 11144
rect 597 11076 729 11110
rect 597 11042 646 11076
rect 680 11042 729 11076
rect 597 11008 729 11042
rect 597 10974 646 11008
rect 680 10974 729 11008
rect 597 10940 729 10974
rect 597 10906 646 10940
rect 680 10906 729 10940
rect 597 10872 729 10906
rect 597 10838 646 10872
rect 680 10838 729 10872
rect 597 10804 729 10838
rect 597 10770 646 10804
rect 680 10770 729 10804
rect 597 10736 729 10770
rect 597 10702 646 10736
rect 680 10702 729 10736
rect 597 10668 729 10702
rect 597 10634 646 10668
rect 680 10634 729 10668
rect 597 10600 729 10634
rect 597 10566 646 10600
rect 680 10566 729 10600
rect 597 10532 729 10566
rect 597 10498 646 10532
rect 680 10498 729 10532
rect 597 10464 729 10498
rect 597 10430 646 10464
rect 680 10430 729 10464
rect 597 10396 729 10430
rect 597 10362 646 10396
rect 680 10362 729 10396
rect 597 10328 729 10362
rect 597 10294 646 10328
rect 680 10294 729 10328
rect 597 10260 729 10294
rect 597 10226 646 10260
rect 680 10226 729 10260
rect 597 10192 729 10226
rect 14247 34672 14381 34706
rect 14247 34638 14297 34672
rect 14331 34638 14381 34672
rect 14247 34604 14381 34638
rect 14247 34570 14297 34604
rect 14331 34570 14381 34604
rect 14247 34536 14381 34570
rect 14247 34502 14297 34536
rect 14331 34502 14381 34536
rect 14247 34468 14381 34502
rect 14247 34434 14297 34468
rect 14331 34434 14381 34468
rect 14247 34400 14381 34434
rect 14247 34366 14297 34400
rect 14331 34366 14381 34400
rect 14247 34332 14381 34366
rect 14247 34298 14297 34332
rect 14331 34298 14381 34332
rect 14247 34264 14381 34298
rect 14247 34230 14297 34264
rect 14331 34230 14381 34264
rect 14247 34196 14381 34230
rect 14247 34162 14297 34196
rect 14331 34162 14381 34196
rect 14247 34128 14381 34162
rect 14247 34094 14297 34128
rect 14331 34094 14381 34128
rect 14247 34060 14381 34094
rect 14247 34026 14297 34060
rect 14331 34026 14381 34060
rect 14247 33992 14381 34026
rect 14247 33958 14297 33992
rect 14331 33958 14381 33992
rect 14247 33924 14381 33958
rect 14247 33890 14297 33924
rect 14331 33890 14381 33924
rect 14247 33856 14381 33890
rect 14247 33822 14297 33856
rect 14331 33822 14381 33856
rect 14247 33788 14381 33822
rect 14247 33754 14297 33788
rect 14331 33754 14381 33788
rect 14247 33720 14381 33754
rect 14247 33686 14297 33720
rect 14331 33686 14381 33720
rect 14247 33652 14381 33686
rect 14247 33618 14297 33652
rect 14331 33618 14381 33652
rect 14247 33584 14381 33618
rect 14247 33550 14297 33584
rect 14331 33550 14381 33584
rect 14247 33516 14381 33550
rect 14247 33482 14297 33516
rect 14331 33482 14381 33516
rect 14247 33448 14381 33482
rect 14247 33414 14297 33448
rect 14331 33414 14381 33448
rect 14247 33380 14381 33414
rect 14247 33346 14297 33380
rect 14331 33346 14381 33380
rect 14247 33312 14381 33346
rect 14247 33278 14297 33312
rect 14331 33278 14381 33312
rect 14247 33244 14381 33278
rect 14247 33210 14297 33244
rect 14331 33210 14381 33244
rect 14247 33176 14381 33210
rect 14247 33142 14297 33176
rect 14331 33142 14381 33176
rect 14247 33108 14381 33142
rect 14247 33074 14297 33108
rect 14331 33074 14381 33108
rect 14247 33040 14381 33074
rect 14247 33006 14297 33040
rect 14331 33006 14381 33040
rect 14247 32972 14381 33006
rect 14247 32938 14297 32972
rect 14331 32938 14381 32972
rect 14247 32904 14381 32938
rect 14247 32870 14297 32904
rect 14331 32870 14381 32904
rect 14247 32836 14381 32870
rect 14247 32802 14297 32836
rect 14331 32802 14381 32836
rect 14247 32768 14381 32802
rect 14247 32734 14297 32768
rect 14331 32734 14381 32768
rect 14247 32700 14381 32734
rect 14247 32666 14297 32700
rect 14331 32666 14381 32700
rect 14247 32632 14381 32666
rect 14247 32598 14297 32632
rect 14331 32598 14381 32632
rect 14247 32564 14381 32598
rect 14247 32530 14297 32564
rect 14331 32530 14381 32564
rect 14247 32496 14381 32530
rect 14247 32462 14297 32496
rect 14331 32462 14381 32496
rect 14247 32428 14381 32462
rect 14247 32394 14297 32428
rect 14331 32394 14381 32428
rect 14247 32360 14381 32394
rect 14247 32326 14297 32360
rect 14331 32326 14381 32360
rect 14247 32292 14381 32326
rect 14247 32258 14297 32292
rect 14331 32258 14381 32292
rect 14247 32224 14381 32258
rect 14247 32190 14297 32224
rect 14331 32190 14381 32224
rect 14247 32156 14381 32190
rect 14247 32122 14297 32156
rect 14331 32122 14381 32156
rect 14247 32088 14381 32122
rect 14247 32054 14297 32088
rect 14331 32054 14381 32088
rect 14247 32020 14381 32054
rect 14247 31986 14297 32020
rect 14331 31986 14381 32020
rect 14247 31952 14381 31986
rect 14247 31918 14297 31952
rect 14331 31918 14381 31952
rect 14247 31884 14381 31918
rect 14247 31850 14297 31884
rect 14331 31850 14381 31884
rect 14247 31816 14381 31850
rect 14247 31782 14297 31816
rect 14331 31782 14381 31816
rect 14247 31748 14381 31782
rect 14247 31714 14297 31748
rect 14331 31714 14381 31748
rect 14247 31680 14381 31714
rect 14247 31646 14297 31680
rect 14331 31646 14381 31680
rect 14247 31612 14381 31646
rect 14247 31578 14297 31612
rect 14331 31578 14381 31612
rect 14247 31544 14381 31578
rect 14247 31510 14297 31544
rect 14331 31510 14381 31544
rect 14247 31476 14381 31510
rect 14247 31442 14297 31476
rect 14331 31442 14381 31476
rect 14247 31408 14381 31442
rect 14247 31374 14297 31408
rect 14331 31374 14381 31408
rect 14247 31340 14381 31374
rect 14247 31306 14297 31340
rect 14331 31306 14381 31340
rect 14247 31272 14381 31306
rect 14247 31238 14297 31272
rect 14331 31238 14381 31272
rect 14247 31204 14381 31238
rect 14247 31170 14297 31204
rect 14331 31170 14381 31204
rect 14247 31136 14381 31170
rect 14247 31102 14297 31136
rect 14331 31102 14381 31136
rect 14247 31068 14381 31102
rect 14247 31034 14297 31068
rect 14331 31034 14381 31068
rect 14247 31000 14381 31034
rect 14247 30966 14297 31000
rect 14331 30966 14381 31000
rect 14247 30932 14381 30966
rect 14247 30898 14297 30932
rect 14331 30898 14381 30932
rect 14247 30864 14381 30898
rect 14247 30830 14297 30864
rect 14331 30830 14381 30864
rect 14247 30796 14381 30830
rect 14247 30762 14297 30796
rect 14331 30762 14381 30796
rect 14247 30728 14381 30762
rect 14247 30694 14297 30728
rect 14331 30694 14381 30728
rect 14247 30660 14381 30694
rect 14247 30626 14297 30660
rect 14331 30626 14381 30660
rect 14247 30592 14381 30626
rect 14247 30558 14297 30592
rect 14331 30558 14381 30592
rect 14247 30524 14381 30558
rect 14247 30490 14297 30524
rect 14331 30490 14381 30524
rect 14247 30456 14381 30490
rect 14247 30422 14297 30456
rect 14331 30422 14381 30456
rect 14247 30388 14381 30422
rect 14247 30354 14297 30388
rect 14331 30354 14381 30388
rect 14247 30320 14381 30354
rect 14247 30286 14297 30320
rect 14331 30286 14381 30320
rect 14247 30252 14381 30286
rect 14247 30218 14297 30252
rect 14331 30218 14381 30252
rect 14247 30184 14381 30218
rect 14247 30150 14297 30184
rect 14331 30150 14381 30184
rect 14247 30116 14381 30150
rect 14247 30082 14297 30116
rect 14331 30082 14381 30116
rect 14247 30048 14381 30082
rect 14247 30014 14297 30048
rect 14331 30014 14381 30048
rect 14247 29980 14381 30014
rect 14247 29946 14297 29980
rect 14331 29946 14381 29980
rect 14247 29912 14381 29946
rect 14247 29878 14297 29912
rect 14331 29878 14381 29912
rect 14247 29844 14381 29878
rect 14247 29810 14297 29844
rect 14331 29810 14381 29844
rect 14247 29776 14381 29810
rect 14247 29742 14297 29776
rect 14331 29742 14381 29776
rect 14247 29708 14381 29742
rect 14247 29674 14297 29708
rect 14331 29674 14381 29708
rect 14247 29640 14381 29674
rect 14247 29606 14297 29640
rect 14331 29606 14381 29640
rect 14247 29572 14381 29606
rect 14247 29538 14297 29572
rect 14331 29538 14381 29572
rect 14247 29504 14381 29538
rect 14247 29470 14297 29504
rect 14331 29470 14381 29504
rect 14247 29436 14381 29470
rect 14247 29402 14297 29436
rect 14331 29402 14381 29436
rect 14247 29368 14381 29402
rect 14247 29334 14297 29368
rect 14331 29334 14381 29368
rect 14247 29300 14381 29334
rect 14247 29266 14297 29300
rect 14331 29266 14381 29300
rect 14247 29232 14381 29266
rect 14247 29198 14297 29232
rect 14331 29198 14381 29232
rect 14247 29164 14381 29198
rect 14247 29130 14297 29164
rect 14331 29130 14381 29164
rect 14247 29096 14381 29130
rect 14247 29062 14297 29096
rect 14331 29062 14381 29096
rect 14247 29028 14381 29062
rect 14247 28994 14297 29028
rect 14331 28994 14381 29028
rect 14247 28960 14381 28994
rect 14247 28926 14297 28960
rect 14331 28926 14381 28960
rect 14247 28892 14381 28926
rect 14247 28858 14297 28892
rect 14331 28858 14381 28892
rect 14247 28824 14381 28858
rect 14247 28790 14297 28824
rect 14331 28790 14381 28824
rect 14247 28756 14381 28790
rect 14247 28722 14297 28756
rect 14331 28722 14381 28756
rect 14247 28688 14381 28722
rect 14247 28654 14297 28688
rect 14331 28654 14381 28688
rect 14247 28620 14381 28654
rect 14247 28586 14297 28620
rect 14331 28586 14381 28620
rect 14247 28552 14381 28586
rect 14247 28518 14297 28552
rect 14331 28518 14381 28552
rect 14247 28484 14381 28518
rect 14247 28450 14297 28484
rect 14331 28450 14381 28484
rect 14247 28416 14381 28450
rect 14247 28382 14297 28416
rect 14331 28382 14381 28416
rect 14247 28348 14381 28382
rect 14247 28314 14297 28348
rect 14331 28314 14381 28348
rect 14247 28280 14381 28314
rect 14247 28246 14297 28280
rect 14331 28246 14381 28280
rect 14247 28212 14381 28246
rect 14247 28178 14297 28212
rect 14331 28178 14381 28212
rect 14247 28144 14381 28178
rect 14247 28110 14297 28144
rect 14331 28110 14381 28144
rect 14247 28076 14381 28110
rect 14247 28042 14297 28076
rect 14331 28042 14381 28076
rect 14247 28008 14381 28042
rect 14247 27974 14297 28008
rect 14331 27974 14381 28008
rect 14247 27940 14381 27974
rect 14247 27906 14297 27940
rect 14331 27906 14381 27940
rect 14247 27872 14381 27906
rect 14247 27838 14297 27872
rect 14331 27838 14381 27872
rect 14247 27804 14381 27838
rect 14247 27770 14297 27804
rect 14331 27770 14381 27804
rect 14247 27736 14381 27770
rect 14247 27702 14297 27736
rect 14331 27702 14381 27736
rect 14247 27668 14381 27702
rect 14247 27634 14297 27668
rect 14331 27634 14381 27668
rect 14247 27600 14381 27634
rect 14247 27566 14297 27600
rect 14331 27566 14381 27600
rect 14247 27532 14381 27566
rect 14247 27498 14297 27532
rect 14331 27498 14381 27532
rect 14247 27464 14381 27498
rect 14247 27430 14297 27464
rect 14331 27430 14381 27464
rect 14247 27396 14381 27430
rect 14247 27362 14297 27396
rect 14331 27362 14381 27396
rect 14247 27328 14381 27362
rect 14247 27294 14297 27328
rect 14331 27294 14381 27328
rect 14247 27260 14381 27294
rect 14247 27226 14297 27260
rect 14331 27226 14381 27260
rect 14247 27192 14381 27226
rect 14247 27158 14297 27192
rect 14331 27158 14381 27192
rect 14247 27124 14381 27158
rect 14247 27090 14297 27124
rect 14331 27090 14381 27124
rect 14247 27056 14381 27090
rect 14247 27022 14297 27056
rect 14331 27022 14381 27056
rect 14247 26988 14381 27022
rect 14247 26954 14297 26988
rect 14331 26954 14381 26988
rect 14247 26920 14381 26954
rect 14247 26886 14297 26920
rect 14331 26886 14381 26920
rect 14247 26852 14381 26886
rect 14247 26818 14297 26852
rect 14331 26818 14381 26852
rect 14247 26784 14381 26818
rect 14247 26750 14297 26784
rect 14331 26750 14381 26784
rect 14247 26716 14381 26750
rect 14247 26682 14297 26716
rect 14331 26682 14381 26716
rect 14247 26648 14381 26682
rect 14247 26614 14297 26648
rect 14331 26614 14381 26648
rect 14247 26580 14381 26614
rect 14247 26546 14297 26580
rect 14331 26546 14381 26580
rect 14247 26512 14381 26546
rect 14247 26478 14297 26512
rect 14331 26478 14381 26512
rect 14247 26444 14381 26478
rect 14247 26410 14297 26444
rect 14331 26410 14381 26444
rect 14247 26376 14381 26410
rect 14247 26342 14297 26376
rect 14331 26342 14381 26376
rect 14247 26308 14381 26342
rect 14247 26274 14297 26308
rect 14331 26274 14381 26308
rect 14247 26240 14381 26274
rect 14247 26206 14297 26240
rect 14331 26206 14381 26240
rect 14247 26172 14381 26206
rect 14247 26138 14297 26172
rect 14331 26138 14381 26172
rect 14247 26104 14381 26138
rect 14247 26070 14297 26104
rect 14331 26070 14381 26104
rect 14247 26036 14381 26070
rect 14247 26002 14297 26036
rect 14331 26002 14381 26036
rect 14247 25968 14381 26002
rect 14247 25934 14297 25968
rect 14331 25934 14381 25968
rect 14247 25900 14381 25934
rect 14247 25866 14297 25900
rect 14331 25866 14381 25900
rect 14247 25832 14381 25866
rect 14247 25798 14297 25832
rect 14331 25798 14381 25832
rect 14247 25764 14381 25798
rect 14247 25730 14297 25764
rect 14331 25730 14381 25764
rect 14247 25696 14381 25730
rect 14247 25662 14297 25696
rect 14331 25662 14381 25696
rect 14247 25628 14381 25662
rect 14247 25594 14297 25628
rect 14331 25594 14381 25628
rect 14247 25560 14381 25594
rect 14247 25526 14297 25560
rect 14331 25526 14381 25560
rect 14247 25492 14381 25526
rect 14247 25458 14297 25492
rect 14331 25458 14381 25492
rect 14247 25424 14381 25458
rect 14247 25390 14297 25424
rect 14331 25390 14381 25424
rect 14247 25356 14381 25390
rect 14247 25322 14297 25356
rect 14331 25322 14381 25356
rect 14247 25288 14381 25322
rect 14247 25254 14297 25288
rect 14331 25254 14381 25288
rect 14247 25220 14381 25254
rect 14247 25186 14297 25220
rect 14331 25186 14381 25220
rect 14247 25152 14381 25186
rect 14247 25118 14297 25152
rect 14331 25118 14381 25152
rect 14247 25084 14381 25118
rect 14247 25050 14297 25084
rect 14331 25050 14381 25084
rect 14247 25016 14381 25050
rect 14247 24982 14297 25016
rect 14331 24982 14381 25016
rect 14247 24948 14381 24982
rect 14247 24914 14297 24948
rect 14331 24914 14381 24948
rect 14247 24880 14381 24914
rect 14247 24846 14297 24880
rect 14331 24846 14381 24880
rect 14247 24812 14381 24846
rect 14247 24778 14297 24812
rect 14331 24778 14381 24812
rect 14247 24744 14381 24778
rect 14247 24710 14297 24744
rect 14331 24710 14381 24744
rect 14247 24676 14381 24710
rect 14247 24642 14297 24676
rect 14331 24642 14381 24676
rect 14247 24608 14381 24642
rect 14247 24574 14297 24608
rect 14331 24574 14381 24608
rect 14247 24540 14381 24574
rect 14247 24506 14297 24540
rect 14331 24506 14381 24540
rect 14247 24472 14381 24506
rect 14247 24438 14297 24472
rect 14331 24438 14381 24472
rect 14247 24404 14381 24438
rect 14247 24370 14297 24404
rect 14331 24370 14381 24404
rect 14247 24336 14381 24370
rect 14247 24302 14297 24336
rect 14331 24302 14381 24336
rect 14247 24268 14381 24302
rect 14247 24234 14297 24268
rect 14331 24234 14381 24268
rect 14247 24200 14381 24234
rect 14247 24166 14297 24200
rect 14331 24166 14381 24200
rect 14247 24132 14381 24166
rect 14247 24098 14297 24132
rect 14331 24098 14381 24132
rect 14247 24064 14381 24098
rect 14247 24030 14297 24064
rect 14331 24030 14381 24064
rect 14247 23996 14381 24030
rect 14247 23962 14297 23996
rect 14331 23962 14381 23996
rect 14247 23928 14381 23962
rect 14247 23894 14297 23928
rect 14331 23894 14381 23928
rect 14247 23860 14381 23894
rect 14247 23826 14297 23860
rect 14331 23826 14381 23860
rect 14247 23792 14381 23826
rect 14247 23758 14297 23792
rect 14331 23758 14381 23792
rect 14247 23724 14381 23758
rect 14247 23690 14297 23724
rect 14331 23690 14381 23724
rect 14247 23656 14381 23690
rect 14247 23622 14297 23656
rect 14331 23622 14381 23656
rect 14247 23588 14381 23622
rect 14247 23554 14297 23588
rect 14331 23554 14381 23588
rect 14247 23520 14381 23554
rect 14247 23486 14297 23520
rect 14331 23486 14381 23520
rect 14247 23452 14381 23486
rect 14247 23418 14297 23452
rect 14331 23418 14381 23452
rect 14247 23384 14381 23418
rect 14247 23350 14297 23384
rect 14331 23350 14381 23384
rect 14247 23316 14381 23350
rect 14247 23282 14297 23316
rect 14331 23282 14381 23316
rect 14247 23248 14381 23282
rect 14247 23214 14297 23248
rect 14331 23214 14381 23248
rect 14247 23180 14381 23214
rect 14247 23146 14297 23180
rect 14331 23146 14381 23180
rect 14247 23112 14381 23146
rect 14247 23078 14297 23112
rect 14331 23078 14381 23112
rect 14247 23044 14381 23078
rect 14247 23010 14297 23044
rect 14331 23010 14381 23044
rect 14247 22976 14381 23010
rect 14247 22942 14297 22976
rect 14331 22942 14381 22976
rect 14247 22908 14381 22942
rect 14247 22874 14297 22908
rect 14331 22874 14381 22908
rect 14247 22840 14381 22874
rect 14247 22806 14297 22840
rect 14331 22806 14381 22840
rect 14247 22772 14381 22806
rect 14247 22738 14297 22772
rect 14331 22738 14381 22772
rect 14247 22704 14381 22738
rect 14247 22670 14297 22704
rect 14331 22670 14381 22704
rect 14247 22636 14381 22670
rect 14247 22602 14297 22636
rect 14331 22602 14381 22636
rect 14247 22568 14381 22602
rect 14247 22534 14297 22568
rect 14331 22534 14381 22568
rect 14247 22500 14381 22534
rect 14247 22466 14297 22500
rect 14331 22466 14381 22500
rect 14247 22432 14381 22466
rect 14247 22398 14297 22432
rect 14331 22398 14381 22432
rect 14247 22364 14381 22398
rect 14247 22330 14297 22364
rect 14331 22330 14381 22364
rect 14247 22296 14381 22330
rect 14247 22262 14297 22296
rect 14331 22262 14381 22296
rect 14247 22228 14381 22262
rect 14247 22194 14297 22228
rect 14331 22194 14381 22228
rect 14247 22160 14381 22194
rect 14247 22126 14297 22160
rect 14331 22126 14381 22160
rect 14247 22092 14381 22126
rect 14247 22058 14297 22092
rect 14331 22058 14381 22092
rect 14247 22024 14381 22058
rect 14247 21990 14297 22024
rect 14331 21990 14381 22024
rect 14247 21956 14381 21990
rect 14247 21922 14297 21956
rect 14331 21922 14381 21956
rect 14247 21888 14381 21922
rect 14247 21854 14297 21888
rect 14331 21854 14381 21888
rect 14247 21820 14381 21854
rect 14247 21786 14297 21820
rect 14331 21786 14381 21820
rect 14247 21752 14381 21786
rect 14247 21718 14297 21752
rect 14331 21718 14381 21752
rect 14247 21684 14381 21718
rect 14247 21650 14297 21684
rect 14331 21650 14381 21684
rect 14247 21616 14381 21650
rect 14247 21582 14297 21616
rect 14331 21582 14381 21616
rect 14247 21548 14381 21582
rect 14247 21514 14297 21548
rect 14331 21514 14381 21548
rect 14247 21480 14381 21514
rect 14247 21446 14297 21480
rect 14331 21446 14381 21480
rect 14247 21412 14381 21446
rect 14247 21378 14297 21412
rect 14331 21378 14381 21412
rect 14247 21344 14381 21378
rect 14247 21310 14297 21344
rect 14331 21310 14381 21344
rect 14247 21276 14381 21310
rect 14247 21242 14297 21276
rect 14331 21242 14381 21276
rect 14247 21208 14381 21242
rect 14247 21174 14297 21208
rect 14331 21174 14381 21208
rect 14247 21140 14381 21174
rect 14247 21106 14297 21140
rect 14331 21106 14381 21140
rect 14247 21072 14381 21106
rect 14247 21038 14297 21072
rect 14331 21038 14381 21072
rect 14247 21004 14381 21038
rect 14247 20970 14297 21004
rect 14331 20970 14381 21004
rect 14247 20936 14381 20970
rect 14247 20902 14297 20936
rect 14331 20902 14381 20936
rect 14247 20868 14381 20902
rect 14247 20834 14297 20868
rect 14331 20834 14381 20868
rect 14247 20800 14381 20834
rect 14247 20766 14297 20800
rect 14331 20766 14381 20800
rect 14247 20732 14381 20766
rect 14247 20698 14297 20732
rect 14331 20698 14381 20732
rect 14247 20664 14381 20698
rect 14247 20630 14297 20664
rect 14331 20630 14381 20664
rect 14247 20596 14381 20630
rect 14247 20562 14297 20596
rect 14331 20562 14381 20596
rect 14247 20528 14381 20562
rect 14247 20494 14297 20528
rect 14331 20494 14381 20528
rect 14247 20460 14381 20494
rect 14247 20426 14297 20460
rect 14331 20426 14381 20460
rect 14247 20392 14381 20426
rect 14247 20358 14297 20392
rect 14331 20358 14381 20392
rect 14247 20324 14381 20358
rect 14247 20290 14297 20324
rect 14331 20290 14381 20324
rect 14247 20256 14381 20290
rect 14247 20222 14297 20256
rect 14331 20222 14381 20256
rect 14247 20188 14381 20222
rect 14247 20154 14297 20188
rect 14331 20154 14381 20188
rect 14247 20120 14381 20154
rect 14247 20086 14297 20120
rect 14331 20086 14381 20120
rect 14247 20052 14381 20086
rect 14247 20018 14297 20052
rect 14331 20018 14381 20052
rect 14247 19984 14381 20018
rect 14247 19950 14297 19984
rect 14331 19950 14381 19984
rect 14247 19916 14381 19950
rect 14247 19882 14297 19916
rect 14331 19882 14381 19916
rect 14247 19848 14381 19882
rect 14247 19814 14297 19848
rect 14331 19814 14381 19848
rect 14247 19780 14381 19814
rect 14247 19746 14297 19780
rect 14331 19746 14381 19780
rect 14247 19712 14381 19746
rect 14247 19678 14297 19712
rect 14331 19678 14381 19712
rect 14247 19644 14381 19678
rect 14247 19610 14297 19644
rect 14331 19610 14381 19644
rect 14247 19576 14381 19610
rect 14247 19542 14297 19576
rect 14331 19542 14381 19576
rect 14247 19508 14381 19542
rect 14247 19474 14297 19508
rect 14331 19474 14381 19508
rect 14247 19440 14381 19474
rect 14247 19406 14297 19440
rect 14331 19406 14381 19440
rect 14247 19372 14381 19406
rect 14247 19338 14297 19372
rect 14331 19338 14381 19372
rect 14247 19304 14381 19338
rect 14247 19270 14297 19304
rect 14331 19270 14381 19304
rect 14247 19236 14381 19270
rect 14247 19202 14297 19236
rect 14331 19202 14381 19236
rect 14247 19168 14381 19202
rect 14247 19134 14297 19168
rect 14331 19134 14381 19168
rect 14247 19100 14381 19134
rect 14247 19066 14297 19100
rect 14331 19066 14381 19100
rect 14247 19032 14381 19066
rect 14247 18998 14297 19032
rect 14331 18998 14381 19032
rect 14247 18964 14381 18998
rect 14247 18930 14297 18964
rect 14331 18930 14381 18964
rect 14247 18896 14381 18930
rect 14247 18862 14297 18896
rect 14331 18862 14381 18896
rect 14247 18828 14381 18862
rect 14247 18794 14297 18828
rect 14331 18794 14381 18828
rect 14247 18760 14381 18794
rect 14247 18726 14297 18760
rect 14331 18726 14381 18760
rect 14247 18692 14381 18726
rect 14247 18658 14297 18692
rect 14331 18658 14381 18692
rect 14247 18624 14381 18658
rect 14247 18590 14297 18624
rect 14331 18590 14381 18624
rect 14247 18556 14381 18590
rect 14247 18522 14297 18556
rect 14331 18522 14381 18556
rect 14247 18488 14381 18522
rect 14247 18454 14297 18488
rect 14331 18454 14381 18488
rect 14247 18420 14381 18454
rect 14247 18386 14297 18420
rect 14331 18386 14381 18420
rect 14247 18352 14381 18386
rect 14247 18318 14297 18352
rect 14331 18318 14381 18352
rect 14247 18284 14381 18318
rect 14247 18250 14297 18284
rect 14331 18250 14381 18284
rect 14247 18216 14381 18250
rect 14247 18182 14297 18216
rect 14331 18182 14381 18216
rect 14247 18148 14381 18182
rect 14247 18114 14297 18148
rect 14331 18114 14381 18148
rect 14247 18080 14381 18114
rect 14247 18046 14297 18080
rect 14331 18046 14381 18080
rect 14247 18012 14381 18046
rect 14247 17978 14297 18012
rect 14331 17978 14381 18012
rect 14247 17944 14381 17978
rect 14247 17910 14297 17944
rect 14331 17910 14381 17944
rect 14247 17876 14381 17910
rect 14247 17842 14297 17876
rect 14331 17842 14381 17876
rect 14247 17808 14381 17842
rect 14247 17774 14297 17808
rect 14331 17774 14381 17808
rect 14247 17740 14381 17774
rect 14247 17706 14297 17740
rect 14331 17706 14381 17740
rect 14247 17672 14381 17706
rect 14247 17638 14297 17672
rect 14331 17638 14381 17672
rect 14247 17604 14381 17638
rect 14247 17570 14297 17604
rect 14331 17570 14381 17604
rect 14247 17536 14381 17570
rect 14247 17502 14297 17536
rect 14331 17502 14381 17536
rect 14247 17468 14381 17502
rect 14247 17434 14297 17468
rect 14331 17434 14381 17468
rect 14247 17400 14381 17434
rect 14247 17366 14297 17400
rect 14331 17366 14381 17400
rect 14247 17332 14381 17366
rect 14247 17298 14297 17332
rect 14331 17298 14381 17332
rect 14247 17264 14381 17298
rect 14247 17230 14297 17264
rect 14331 17230 14381 17264
rect 14247 17196 14381 17230
rect 14247 17162 14297 17196
rect 14331 17162 14381 17196
rect 14247 17128 14381 17162
rect 14247 17094 14297 17128
rect 14331 17094 14381 17128
rect 14247 17060 14381 17094
rect 14247 17026 14297 17060
rect 14331 17026 14381 17060
rect 14247 16992 14381 17026
rect 14247 16958 14297 16992
rect 14331 16958 14381 16992
rect 14247 16924 14381 16958
rect 14247 16890 14297 16924
rect 14331 16890 14381 16924
rect 14247 16856 14381 16890
rect 14247 16822 14297 16856
rect 14331 16822 14381 16856
rect 14247 16788 14381 16822
rect 14247 16754 14297 16788
rect 14331 16754 14381 16788
rect 14247 16720 14381 16754
rect 14247 16686 14297 16720
rect 14331 16686 14381 16720
rect 14247 16652 14381 16686
rect 14247 16618 14297 16652
rect 14331 16618 14381 16652
rect 14247 16584 14381 16618
rect 14247 16550 14297 16584
rect 14331 16550 14381 16584
rect 14247 16516 14381 16550
rect 14247 16482 14297 16516
rect 14331 16482 14381 16516
rect 14247 16448 14381 16482
rect 14247 16414 14297 16448
rect 14331 16414 14381 16448
rect 14247 16380 14381 16414
rect 14247 16346 14297 16380
rect 14331 16346 14381 16380
rect 14247 16312 14381 16346
rect 14247 16278 14297 16312
rect 14331 16278 14381 16312
rect 14247 16244 14381 16278
rect 14247 16210 14297 16244
rect 14331 16210 14381 16244
rect 14247 16176 14381 16210
rect 14247 16142 14297 16176
rect 14331 16142 14381 16176
rect 14247 16108 14381 16142
rect 14247 16074 14297 16108
rect 14331 16074 14381 16108
rect 14247 16040 14381 16074
rect 14247 16006 14297 16040
rect 14331 16006 14381 16040
rect 14247 15972 14381 16006
rect 14247 15938 14297 15972
rect 14331 15938 14381 15972
rect 14247 15904 14381 15938
rect 14247 15870 14297 15904
rect 14331 15870 14381 15904
rect 14247 15836 14381 15870
rect 14247 15802 14297 15836
rect 14331 15802 14381 15836
rect 14247 15768 14381 15802
rect 14247 15734 14297 15768
rect 14331 15734 14381 15768
rect 14247 15700 14381 15734
rect 14247 15666 14297 15700
rect 14331 15666 14381 15700
rect 14247 15632 14381 15666
rect 14247 15598 14297 15632
rect 14331 15598 14381 15632
rect 14247 15564 14381 15598
rect 14247 15530 14297 15564
rect 14331 15530 14381 15564
rect 14247 15496 14381 15530
rect 14247 15462 14297 15496
rect 14331 15462 14381 15496
rect 14247 15428 14381 15462
rect 14247 15394 14297 15428
rect 14331 15394 14381 15428
rect 14247 15360 14381 15394
rect 14247 15326 14297 15360
rect 14331 15326 14381 15360
rect 14247 15292 14381 15326
rect 14247 15258 14297 15292
rect 14331 15258 14381 15292
rect 14247 15224 14381 15258
rect 14247 15190 14297 15224
rect 14331 15190 14381 15224
rect 14247 15156 14381 15190
rect 14247 15122 14297 15156
rect 14331 15122 14381 15156
rect 14247 15088 14381 15122
rect 14247 15054 14297 15088
rect 14331 15054 14381 15088
rect 14247 15020 14381 15054
rect 14247 14986 14297 15020
rect 14331 14986 14381 15020
rect 14247 14952 14381 14986
rect 14247 14918 14297 14952
rect 14331 14918 14381 14952
rect 14247 14884 14381 14918
rect 14247 14850 14297 14884
rect 14331 14850 14381 14884
rect 14247 14816 14381 14850
rect 14247 14782 14297 14816
rect 14331 14782 14381 14816
rect 14247 14748 14381 14782
rect 14247 14714 14297 14748
rect 14331 14714 14381 14748
rect 14247 14680 14381 14714
rect 14247 14646 14297 14680
rect 14331 14646 14381 14680
rect 14247 14612 14381 14646
rect 14247 14578 14297 14612
rect 14331 14578 14381 14612
rect 14247 14544 14381 14578
rect 14247 14510 14297 14544
rect 14331 14510 14381 14544
rect 14247 14476 14381 14510
rect 14247 14442 14297 14476
rect 14331 14442 14381 14476
rect 14247 14408 14381 14442
rect 14247 14374 14297 14408
rect 14331 14374 14381 14408
rect 14247 14340 14381 14374
rect 14247 14306 14297 14340
rect 14331 14306 14381 14340
rect 14247 14272 14381 14306
rect 14247 14238 14297 14272
rect 14331 14238 14381 14272
rect 14247 14204 14381 14238
rect 14247 14170 14297 14204
rect 14331 14170 14381 14204
rect 14247 14136 14381 14170
rect 14247 14102 14297 14136
rect 14331 14102 14381 14136
rect 14247 14068 14381 14102
rect 14247 14034 14297 14068
rect 14331 14034 14381 14068
rect 14247 14000 14381 14034
rect 14247 13966 14297 14000
rect 14331 13966 14381 14000
rect 14247 13932 14381 13966
rect 14247 13898 14297 13932
rect 14331 13898 14381 13932
rect 14247 13864 14381 13898
rect 14247 13830 14297 13864
rect 14331 13830 14381 13864
rect 14247 13796 14381 13830
rect 14247 13762 14297 13796
rect 14331 13762 14381 13796
rect 14247 13728 14381 13762
rect 14247 13694 14297 13728
rect 14331 13694 14381 13728
rect 14247 13660 14381 13694
rect 14247 13626 14297 13660
rect 14331 13626 14381 13660
rect 14247 13592 14381 13626
rect 14247 13558 14297 13592
rect 14331 13558 14381 13592
rect 14247 13524 14381 13558
rect 14247 13490 14297 13524
rect 14331 13490 14381 13524
rect 14247 13456 14381 13490
rect 14247 13422 14297 13456
rect 14331 13422 14381 13456
rect 14247 13388 14381 13422
rect 14247 13354 14297 13388
rect 14331 13354 14381 13388
rect 14247 13320 14381 13354
rect 14247 13286 14297 13320
rect 14331 13286 14381 13320
rect 14247 13252 14381 13286
rect 14247 13218 14297 13252
rect 14331 13218 14381 13252
rect 14247 13184 14381 13218
rect 14247 13150 14297 13184
rect 14331 13150 14381 13184
rect 14247 13116 14381 13150
rect 14247 13082 14297 13116
rect 14331 13082 14381 13116
rect 14247 13048 14381 13082
rect 14247 13014 14297 13048
rect 14331 13014 14381 13048
rect 14247 12980 14381 13014
rect 14247 12946 14297 12980
rect 14331 12946 14381 12980
rect 14247 12912 14381 12946
rect 14247 12878 14297 12912
rect 14331 12878 14381 12912
rect 14247 12844 14381 12878
rect 14247 12810 14297 12844
rect 14331 12810 14381 12844
rect 14247 12776 14381 12810
rect 14247 12742 14297 12776
rect 14331 12742 14381 12776
rect 14247 12708 14381 12742
rect 14247 12674 14297 12708
rect 14331 12674 14381 12708
rect 14247 12640 14381 12674
rect 14247 12606 14297 12640
rect 14331 12606 14381 12640
rect 14247 12572 14381 12606
rect 14247 12538 14297 12572
rect 14331 12538 14381 12572
rect 14247 12504 14381 12538
rect 14247 12470 14297 12504
rect 14331 12470 14381 12504
rect 14247 12436 14381 12470
rect 14247 12402 14297 12436
rect 14331 12402 14381 12436
rect 14247 12368 14381 12402
rect 14247 12334 14297 12368
rect 14331 12334 14381 12368
rect 14247 12300 14381 12334
rect 14247 12266 14297 12300
rect 14331 12266 14381 12300
rect 14247 12232 14381 12266
rect 14247 12198 14297 12232
rect 14331 12198 14381 12232
rect 14247 12164 14381 12198
rect 14247 12130 14297 12164
rect 14331 12130 14381 12164
rect 14247 12096 14381 12130
rect 14247 12062 14297 12096
rect 14331 12062 14381 12096
rect 14247 12028 14381 12062
rect 14247 11994 14297 12028
rect 14331 11994 14381 12028
rect 14247 11960 14381 11994
rect 14247 11926 14297 11960
rect 14331 11926 14381 11960
rect 14247 11892 14381 11926
rect 14247 11858 14297 11892
rect 14331 11858 14381 11892
rect 14247 11824 14381 11858
rect 14247 11790 14297 11824
rect 14331 11790 14381 11824
rect 14247 11756 14381 11790
rect 14247 11722 14297 11756
rect 14331 11722 14381 11756
rect 14247 11688 14381 11722
rect 14247 11654 14297 11688
rect 14331 11654 14381 11688
rect 14247 11620 14381 11654
rect 14247 11586 14297 11620
rect 14331 11586 14381 11620
rect 14247 11552 14381 11586
rect 14247 11518 14297 11552
rect 14331 11518 14381 11552
rect 14247 11484 14381 11518
rect 14247 11450 14297 11484
rect 14331 11450 14381 11484
rect 14247 11416 14381 11450
rect 14247 11382 14297 11416
rect 14331 11382 14381 11416
rect 14247 11348 14381 11382
rect 14247 11314 14297 11348
rect 14331 11314 14381 11348
rect 14247 11280 14381 11314
rect 14247 11246 14297 11280
rect 14331 11246 14381 11280
rect 14247 11212 14381 11246
rect 14247 11178 14297 11212
rect 14331 11178 14381 11212
rect 14247 11144 14381 11178
rect 14247 11110 14297 11144
rect 14331 11110 14381 11144
rect 14247 11076 14381 11110
rect 14247 11042 14297 11076
rect 14331 11042 14381 11076
rect 14247 11008 14381 11042
rect 14247 10974 14297 11008
rect 14331 10974 14381 11008
rect 14247 10940 14381 10974
rect 14247 10906 14297 10940
rect 14331 10906 14381 10940
rect 14247 10872 14381 10906
rect 14247 10838 14297 10872
rect 14331 10838 14381 10872
rect 14247 10804 14381 10838
rect 14247 10770 14297 10804
rect 14331 10770 14381 10804
rect 14247 10736 14381 10770
rect 14247 10702 14297 10736
rect 14331 10702 14381 10736
rect 14247 10668 14381 10702
rect 14247 10634 14297 10668
rect 14331 10634 14381 10668
rect 14247 10600 14381 10634
rect 14247 10566 14297 10600
rect 14331 10566 14381 10600
rect 14247 10532 14381 10566
rect 14247 10498 14297 10532
rect 14331 10498 14381 10532
rect 14247 10464 14381 10498
rect 14247 10430 14297 10464
rect 14331 10430 14381 10464
rect 14247 10396 14381 10430
rect 14247 10362 14297 10396
rect 14331 10362 14381 10396
rect 14247 10328 14381 10362
rect 14247 10294 14297 10328
rect 14331 10294 14381 10328
rect 14247 10260 14381 10294
rect 14247 10226 14297 10260
rect 14331 10226 14381 10260
rect 597 10158 646 10192
rect 680 10158 729 10192
rect 597 10124 729 10158
rect 597 10090 646 10124
rect 680 10090 729 10124
rect 597 10056 729 10090
rect 597 10022 646 10056
rect 680 10022 729 10056
rect 597 9988 729 10022
rect 597 9954 646 9988
rect 680 9954 729 9988
rect 597 9920 729 9954
rect 597 9886 646 9920
rect 680 9886 729 9920
rect 597 9825 729 9886
rect 14247 10192 14381 10226
rect 14247 10158 14297 10192
rect 14331 10158 14381 10192
rect 14247 10124 14381 10158
rect 14247 10090 14297 10124
rect 14331 10090 14381 10124
rect 14247 10056 14381 10090
rect 14247 10022 14297 10056
rect 14331 10022 14381 10056
rect 14247 9988 14381 10022
rect 14247 9954 14297 9988
rect 14331 9954 14381 9988
rect 14247 9920 14381 9954
rect 14247 9886 14297 9920
rect 14331 9886 14381 9920
rect 14247 9825 14381 9886
rect 597 9775 14381 9825
rect 597 9741 773 9775
rect 807 9741 841 9775
rect 875 9741 909 9775
rect 943 9741 977 9775
rect 1011 9741 1045 9775
rect 1079 9741 1113 9775
rect 1147 9741 1181 9775
rect 1215 9741 1249 9775
rect 1283 9741 1317 9775
rect 1351 9741 1385 9775
rect 1419 9741 1453 9775
rect 1487 9741 1521 9775
rect 1555 9741 1589 9775
rect 1623 9741 1657 9775
rect 1691 9741 1725 9775
rect 1759 9741 1793 9775
rect 1827 9741 1861 9775
rect 1895 9741 1929 9775
rect 1963 9741 1997 9775
rect 2031 9741 2065 9775
rect 2099 9741 2133 9775
rect 2167 9741 2201 9775
rect 2235 9741 2269 9775
rect 2303 9741 2337 9775
rect 2371 9741 2405 9775
rect 2439 9741 2473 9775
rect 2507 9741 2541 9775
rect 2575 9741 2609 9775
rect 2643 9741 2677 9775
rect 2711 9741 2745 9775
rect 2779 9741 2813 9775
rect 2847 9741 2881 9775
rect 2915 9741 2949 9775
rect 2983 9741 3017 9775
rect 3051 9741 3085 9775
rect 3119 9741 3153 9775
rect 3187 9741 3221 9775
rect 3255 9741 3289 9775
rect 3323 9741 3357 9775
rect 3391 9741 3425 9775
rect 3459 9741 3493 9775
rect 3527 9741 3561 9775
rect 3595 9741 3629 9775
rect 3663 9741 3697 9775
rect 3731 9741 3765 9775
rect 3799 9741 3833 9775
rect 3867 9741 3901 9775
rect 3935 9741 3969 9775
rect 4003 9741 4037 9775
rect 4071 9741 4105 9775
rect 4139 9741 4173 9775
rect 4207 9741 4241 9775
rect 4275 9741 4309 9775
rect 4343 9741 4377 9775
rect 4411 9741 4445 9775
rect 4479 9741 4513 9775
rect 4547 9741 4581 9775
rect 4615 9741 4649 9775
rect 4683 9741 4717 9775
rect 4751 9741 4785 9775
rect 4819 9741 4853 9775
rect 4887 9741 4921 9775
rect 4955 9741 4989 9775
rect 5023 9741 5057 9775
rect 5091 9741 5125 9775
rect 5159 9741 5193 9775
rect 5227 9741 5261 9775
rect 5295 9741 5329 9775
rect 5363 9741 5397 9775
rect 5431 9741 5465 9775
rect 5499 9741 5533 9775
rect 5567 9741 5601 9775
rect 5635 9741 5669 9775
rect 5703 9741 5737 9775
rect 5771 9741 5805 9775
rect 5839 9741 5873 9775
rect 5907 9741 5941 9775
rect 5975 9741 6009 9775
rect 6043 9741 6077 9775
rect 6111 9741 6145 9775
rect 6179 9741 6213 9775
rect 6247 9741 6281 9775
rect 6315 9741 6349 9775
rect 6383 9741 6417 9775
rect 6451 9741 6485 9775
rect 6519 9741 6553 9775
rect 6587 9741 6621 9775
rect 6655 9741 6689 9775
rect 6723 9741 6757 9775
rect 6791 9741 6825 9775
rect 6859 9741 6893 9775
rect 6927 9741 6961 9775
rect 6995 9741 7029 9775
rect 7063 9741 7097 9775
rect 7131 9741 7165 9775
rect 7199 9741 7233 9775
rect 7267 9741 7301 9775
rect 7335 9741 7369 9775
rect 7403 9741 7437 9775
rect 7471 9741 7505 9775
rect 7539 9741 7573 9775
rect 7607 9741 7641 9775
rect 7675 9741 7709 9775
rect 7743 9741 7777 9775
rect 7811 9741 7845 9775
rect 7879 9741 7913 9775
rect 7947 9741 7981 9775
rect 8015 9741 8049 9775
rect 8083 9741 8117 9775
rect 8151 9741 8185 9775
rect 8219 9741 8253 9775
rect 8287 9741 8321 9775
rect 8355 9741 8389 9775
rect 8423 9741 8457 9775
rect 8491 9741 8525 9775
rect 8559 9741 8593 9775
rect 8627 9741 8661 9775
rect 8695 9741 8729 9775
rect 8763 9741 8797 9775
rect 8831 9741 8865 9775
rect 8899 9741 8933 9775
rect 8967 9741 9001 9775
rect 9035 9741 9069 9775
rect 9103 9741 9137 9775
rect 9171 9741 9205 9775
rect 9239 9741 9273 9775
rect 9307 9741 9341 9775
rect 9375 9741 9409 9775
rect 9443 9741 9477 9775
rect 9511 9741 9545 9775
rect 9579 9741 9613 9775
rect 9647 9741 9681 9775
rect 9715 9741 9749 9775
rect 9783 9741 9817 9775
rect 9851 9741 9885 9775
rect 9919 9741 9953 9775
rect 9987 9741 10021 9775
rect 10055 9741 10089 9775
rect 10123 9741 10157 9775
rect 10191 9741 10225 9775
rect 10259 9741 10293 9775
rect 10327 9741 10361 9775
rect 10395 9741 10429 9775
rect 10463 9741 10497 9775
rect 10531 9741 10565 9775
rect 10599 9741 10633 9775
rect 10667 9741 10701 9775
rect 10735 9741 10769 9775
rect 10803 9741 10837 9775
rect 10871 9741 10905 9775
rect 10939 9741 10973 9775
rect 11007 9741 11041 9775
rect 11075 9741 11109 9775
rect 11143 9741 11177 9775
rect 11211 9741 11245 9775
rect 11279 9741 11313 9775
rect 11347 9741 11381 9775
rect 11415 9741 11449 9775
rect 11483 9741 11517 9775
rect 11551 9741 11585 9775
rect 11619 9741 11653 9775
rect 11687 9741 11721 9775
rect 11755 9741 11789 9775
rect 11823 9741 11857 9775
rect 11891 9741 11925 9775
rect 11959 9741 11993 9775
rect 12027 9741 12061 9775
rect 12095 9741 12129 9775
rect 12163 9741 12197 9775
rect 12231 9741 12265 9775
rect 12299 9741 12333 9775
rect 12367 9741 12401 9775
rect 12435 9741 12469 9775
rect 12503 9741 12537 9775
rect 12571 9741 12605 9775
rect 12639 9741 12673 9775
rect 12707 9741 12741 9775
rect 12775 9741 12809 9775
rect 12843 9741 12877 9775
rect 12911 9741 12945 9775
rect 12979 9741 13013 9775
rect 13047 9741 13081 9775
rect 13115 9741 13149 9775
rect 13183 9741 13217 9775
rect 13251 9741 13285 9775
rect 13319 9741 13353 9775
rect 13387 9741 13421 9775
rect 13455 9741 13489 9775
rect 13523 9741 13557 9775
rect 13591 9741 13625 9775
rect 13659 9741 13693 9775
rect 13727 9741 13761 9775
rect 13795 9741 13829 9775
rect 13863 9741 13897 9775
rect 13931 9741 13965 9775
rect 13999 9741 14033 9775
rect 14067 9741 14101 9775
rect 14135 9741 14169 9775
rect 14203 9741 14381 9775
rect 597 9691 14381 9741
<< mvpsubdiffcont >>
rect 492 36465 526 36499
rect 560 36465 594 36499
rect 628 36465 662 36499
rect 696 36465 730 36499
rect 764 36465 798 36499
rect 832 36465 866 36499
rect 900 36465 934 36499
rect 968 36465 1002 36499
rect 1036 36465 1070 36499
rect 1104 36465 1138 36499
rect 1172 36465 1206 36499
rect 1240 36465 1274 36499
rect 1308 36465 1342 36499
rect 1376 36465 1410 36499
rect 1444 36465 1478 36499
rect 1512 36465 1546 36499
rect 1580 36465 1614 36499
rect 1648 36465 1682 36499
rect 1716 36465 1750 36499
rect 1784 36465 1818 36499
rect 1852 36465 1886 36499
rect 1920 36465 1954 36499
rect 1988 36465 2022 36499
rect 2056 36465 2090 36499
rect 2124 36465 2158 36499
rect 2192 36465 2226 36499
rect 2260 36465 2294 36499
rect 2328 36465 2362 36499
rect 2396 36465 2430 36499
rect 2464 36465 2498 36499
rect 2532 36465 2566 36499
rect 2600 36465 2634 36499
rect 2668 36465 2702 36499
rect 2736 36465 2770 36499
rect 2804 36465 2838 36499
rect 2872 36465 2906 36499
rect 2940 36465 2974 36499
rect 3008 36465 3042 36499
rect 3076 36465 3110 36499
rect 3144 36465 3178 36499
rect 3212 36465 3246 36499
rect 3280 36465 3314 36499
rect 3348 36465 3382 36499
rect 3416 36465 3450 36499
rect 3484 36465 3518 36499
rect 3552 36465 3586 36499
rect 3620 36465 3654 36499
rect 3688 36465 3722 36499
rect 3756 36465 3790 36499
rect 3824 36465 3858 36499
rect 3892 36465 3926 36499
rect 3960 36465 3994 36499
rect 4028 36465 4062 36499
rect 4096 36465 4130 36499
rect 4164 36465 4198 36499
rect 4232 36465 4266 36499
rect 4300 36465 4334 36499
rect 4368 36465 4402 36499
rect 4436 36465 4470 36499
rect 4504 36465 4538 36499
rect 4572 36465 4606 36499
rect 4640 36465 4674 36499
rect 4708 36465 4742 36499
rect 4776 36465 4810 36499
rect 4844 36465 4878 36499
rect 4912 36465 4946 36499
rect 4980 36465 5014 36499
rect 5048 36465 5082 36499
rect 5116 36465 5150 36499
rect 5184 36465 5218 36499
rect 5252 36465 5286 36499
rect 5320 36465 5354 36499
rect 5388 36465 5422 36499
rect 5456 36465 5490 36499
rect 5524 36465 5558 36499
rect 5592 36465 5626 36499
rect 5660 36465 5694 36499
rect 5728 36465 5762 36499
rect 5796 36465 5830 36499
rect 5864 36465 5898 36499
rect 5932 36465 5966 36499
rect 6000 36465 6034 36499
rect 6068 36465 6102 36499
rect 6136 36465 6170 36499
rect 6204 36465 6238 36499
rect 6272 36465 6306 36499
rect 6340 36465 6374 36499
rect 6408 36465 6442 36499
rect 6476 36465 6510 36499
rect 6544 36465 6578 36499
rect 6612 36465 6646 36499
rect 6680 36465 6714 36499
rect 6748 36465 6782 36499
rect 6816 36465 6850 36499
rect 6884 36465 6918 36499
rect 6952 36465 6986 36499
rect 7020 36465 7054 36499
rect 7088 36465 7122 36499
rect 7156 36465 7190 36499
rect 7224 36465 7258 36499
rect 7292 36465 7326 36499
rect 7360 36465 7394 36499
rect 7428 36465 7462 36499
rect 7496 36465 7530 36499
rect 7564 36465 7598 36499
rect 7632 36465 7666 36499
rect 7700 36465 7734 36499
rect 7768 36465 7802 36499
rect 7836 36465 7870 36499
rect 7904 36465 7938 36499
rect 7972 36465 8006 36499
rect 8040 36465 8074 36499
rect 8108 36465 8142 36499
rect 8176 36465 8210 36499
rect 8244 36465 8278 36499
rect 8312 36465 8346 36499
rect 8380 36465 8414 36499
rect 8448 36465 8482 36499
rect 8516 36465 8550 36499
rect 8584 36465 8618 36499
rect 8652 36465 8686 36499
rect 8720 36465 8754 36499
rect 8788 36465 8822 36499
rect 8856 36465 8890 36499
rect 8924 36465 8958 36499
rect 8992 36465 9026 36499
rect 9060 36465 9094 36499
rect 9128 36465 9162 36499
rect 9196 36465 9230 36499
rect 9264 36465 9298 36499
rect 9332 36465 9366 36499
rect 9400 36465 9434 36499
rect 9468 36465 9502 36499
rect 9536 36465 9570 36499
rect 9604 36465 9638 36499
rect 9672 36465 9706 36499
rect 9740 36465 9774 36499
rect 9808 36465 9842 36499
rect 9876 36465 9910 36499
rect 9944 36465 9978 36499
rect 10012 36465 10046 36499
rect 10080 36465 10114 36499
rect 10148 36465 10182 36499
rect 10216 36465 10250 36499
rect 10284 36465 10318 36499
rect 10352 36465 10386 36499
rect 10420 36465 10454 36499
rect 10488 36465 10522 36499
rect 10556 36465 10590 36499
rect 10624 36465 10658 36499
rect 10692 36465 10726 36499
rect 10760 36465 10794 36499
rect 10828 36465 10862 36499
rect 10896 36465 10930 36499
rect 10964 36465 10998 36499
rect 11032 36465 11066 36499
rect 11100 36465 11134 36499
rect 11168 36465 11202 36499
rect 11236 36465 11270 36499
rect 11304 36465 11338 36499
rect 11372 36465 11406 36499
rect 11440 36465 11474 36499
rect 11508 36465 11542 36499
rect 11576 36465 11610 36499
rect 11644 36465 11678 36499
rect 11712 36465 11746 36499
rect 11780 36465 11814 36499
rect 11848 36465 11882 36499
rect 11916 36465 11950 36499
rect 11984 36465 12018 36499
rect 12052 36465 12086 36499
rect 12120 36465 12154 36499
rect 12188 36465 12222 36499
rect 12256 36465 12290 36499
rect 12324 36465 12358 36499
rect 12392 36465 12426 36499
rect 12460 36465 12494 36499
rect 12528 36465 12562 36499
rect 12596 36465 12630 36499
rect 12664 36465 12698 36499
rect 12732 36465 12766 36499
rect 12800 36465 12834 36499
rect 12868 36465 12902 36499
rect 12936 36465 12970 36499
rect 13004 36465 13038 36499
rect 13072 36465 13106 36499
rect 13140 36465 13174 36499
rect 13208 36465 13242 36499
rect 13276 36465 13310 36499
rect 13344 36465 13378 36499
rect 13412 36465 13446 36499
rect 13480 36465 13514 36499
rect 13548 36465 13582 36499
rect 13616 36465 13650 36499
rect 13684 36465 13718 36499
rect 13752 36465 13786 36499
rect 13820 36465 13854 36499
rect 13888 36465 13922 36499
rect 13956 36465 13990 36499
rect 14024 36465 14058 36499
rect 14092 36465 14126 36499
rect 14160 36465 14194 36499
rect 14228 36465 14262 36499
rect 14296 36465 14330 36499
rect 14364 36465 14398 36499
rect 14432 36465 14466 36499
rect 322 36301 356 36335
rect 322 36233 356 36267
rect 14609 36293 14643 36327
rect 322 36165 356 36199
rect 322 36097 356 36131
rect 322 36029 356 36063
rect 322 35961 356 35995
rect 322 35893 356 35927
rect 322 35825 356 35859
rect 322 35757 356 35791
rect 322 35689 356 35723
rect 322 35621 356 35655
rect 322 35553 356 35587
rect 322 35485 356 35519
rect 322 35417 356 35451
rect 322 35349 356 35383
rect 322 35281 356 35315
rect 322 35213 356 35247
rect 322 35145 356 35179
rect 322 35077 356 35111
rect 322 35009 356 35043
rect 322 34941 356 34975
rect 322 34873 356 34907
rect 322 34805 356 34839
rect 322 34737 356 34771
rect 322 34669 356 34703
rect 322 34601 356 34635
rect 322 34533 356 34567
rect 322 34465 356 34499
rect 322 34397 356 34431
rect 322 34329 356 34363
rect 322 34261 356 34295
rect 322 34193 356 34227
rect 322 34125 356 34159
rect 322 34057 356 34091
rect 322 33989 356 34023
rect 322 33921 356 33955
rect 322 33853 356 33887
rect 322 33785 356 33819
rect 322 33717 356 33751
rect 322 33649 356 33683
rect 322 33581 356 33615
rect 322 33513 356 33547
rect 322 33445 356 33479
rect 322 33377 356 33411
rect 322 33309 356 33343
rect 322 33241 356 33275
rect 322 33173 356 33207
rect 322 33105 356 33139
rect 322 33037 356 33071
rect 322 32969 356 33003
rect 322 32901 356 32935
rect 322 32833 356 32867
rect 322 32765 356 32799
rect 322 32697 356 32731
rect 322 32629 356 32663
rect 322 32561 356 32595
rect 322 32493 356 32527
rect 322 32425 356 32459
rect 322 32357 356 32391
rect 322 32289 356 32323
rect 322 32221 356 32255
rect 322 32153 356 32187
rect 322 32085 356 32119
rect 322 32017 356 32051
rect 322 31949 356 31983
rect 322 31881 356 31915
rect 322 31813 356 31847
rect 322 31745 356 31779
rect 322 31677 356 31711
rect 322 31609 356 31643
rect 322 31541 356 31575
rect 322 31473 356 31507
rect 322 31405 356 31439
rect 322 31337 356 31371
rect 322 31269 356 31303
rect 322 31201 356 31235
rect 322 31133 356 31167
rect 322 31065 356 31099
rect 322 30997 356 31031
rect 322 30929 356 30963
rect 322 30861 356 30895
rect 322 30793 356 30827
rect 322 30725 356 30759
rect 322 30657 356 30691
rect 322 30589 356 30623
rect 322 30521 356 30555
rect 322 30453 356 30487
rect 322 30385 356 30419
rect 322 30317 356 30351
rect 322 30249 356 30283
rect 322 30181 356 30215
rect 322 30113 356 30147
rect 322 30045 356 30079
rect 322 29977 356 30011
rect 322 29909 356 29943
rect 322 29841 356 29875
rect 322 29773 356 29807
rect 322 29705 356 29739
rect 322 29637 356 29671
rect 322 29569 356 29603
rect 322 29501 356 29535
rect 322 29433 356 29467
rect 322 29365 356 29399
rect 322 29297 356 29331
rect 322 29229 356 29263
rect 322 29161 356 29195
rect 322 29093 356 29127
rect 322 29025 356 29059
rect 322 28957 356 28991
rect 322 28889 356 28923
rect 322 28821 356 28855
rect 322 28753 356 28787
rect 322 28685 356 28719
rect 322 28617 356 28651
rect 322 28549 356 28583
rect 322 28481 356 28515
rect 322 28413 356 28447
rect 322 28345 356 28379
rect 322 28277 356 28311
rect 322 28209 356 28243
rect 322 28141 356 28175
rect 322 28073 356 28107
rect 322 28005 356 28039
rect 322 27937 356 27971
rect 322 27869 356 27903
rect 322 27801 356 27835
rect 322 27733 356 27767
rect 322 27665 356 27699
rect 322 27597 356 27631
rect 322 27529 356 27563
rect 322 27461 356 27495
rect 322 27393 356 27427
rect 322 27325 356 27359
rect 322 27257 356 27291
rect 322 27189 356 27223
rect 322 27121 356 27155
rect 322 27053 356 27087
rect 322 26985 356 27019
rect 322 26917 356 26951
rect 322 26849 356 26883
rect 322 26781 356 26815
rect 322 26713 356 26747
rect 322 26645 356 26679
rect 322 26577 356 26611
rect 322 26509 356 26543
rect 322 26441 356 26475
rect 322 26373 356 26407
rect 322 26305 356 26339
rect 322 26237 356 26271
rect 322 26169 356 26203
rect 322 26101 356 26135
rect 322 26033 356 26067
rect 322 25965 356 25999
rect 322 25897 356 25931
rect 322 25829 356 25863
rect 322 25761 356 25795
rect 322 25693 356 25727
rect 322 25625 356 25659
rect 322 25557 356 25591
rect 322 25489 356 25523
rect 322 25421 356 25455
rect 322 25353 356 25387
rect 322 25285 356 25319
rect 322 25217 356 25251
rect 322 25149 356 25183
rect 322 25081 356 25115
rect 322 25013 356 25047
rect 322 24945 356 24979
rect 322 24877 356 24911
rect 322 24809 356 24843
rect 322 24741 356 24775
rect 322 24673 356 24707
rect 322 24605 356 24639
rect 322 24537 356 24571
rect 322 24469 356 24503
rect 322 24401 356 24435
rect 322 24333 356 24367
rect 322 24265 356 24299
rect 322 24197 356 24231
rect 322 24129 356 24163
rect 322 24061 356 24095
rect 322 23993 356 24027
rect 322 23925 356 23959
rect 322 23857 356 23891
rect 322 23789 356 23823
rect 322 23721 356 23755
rect 322 23653 356 23687
rect 322 23585 356 23619
rect 322 23517 356 23551
rect 322 23449 356 23483
rect 322 23381 356 23415
rect 322 23313 356 23347
rect 322 23245 356 23279
rect 322 23177 356 23211
rect 322 23109 356 23143
rect 322 23041 356 23075
rect 322 22973 356 23007
rect 322 22905 356 22939
rect 322 22837 356 22871
rect 322 22769 356 22803
rect 322 22701 356 22735
rect 322 22633 356 22667
rect 322 22565 356 22599
rect 322 22497 356 22531
rect 322 22429 356 22463
rect 322 22361 356 22395
rect 322 22293 356 22327
rect 322 22225 356 22259
rect 322 22157 356 22191
rect 322 22089 356 22123
rect 322 22021 356 22055
rect 322 21953 356 21987
rect 322 21885 356 21919
rect 322 21817 356 21851
rect 322 21749 356 21783
rect 322 21681 356 21715
rect 322 21613 356 21647
rect 322 21545 356 21579
rect 322 21477 356 21511
rect 322 21409 356 21443
rect 322 21341 356 21375
rect 322 21273 356 21307
rect 322 21205 356 21239
rect 322 21137 356 21171
rect 322 21069 356 21103
rect 322 21001 356 21035
rect 322 20933 356 20967
rect 322 20865 356 20899
rect 322 20797 356 20831
rect 322 20729 356 20763
rect 322 20661 356 20695
rect 322 20593 356 20627
rect 322 20525 356 20559
rect 322 20457 356 20491
rect 322 20389 356 20423
rect 322 20321 356 20355
rect 322 20253 356 20287
rect 322 20185 356 20219
rect 322 20117 356 20151
rect 322 20049 356 20083
rect 322 19981 356 20015
rect 322 19913 356 19947
rect 322 19845 356 19879
rect 322 19777 356 19811
rect 322 19709 356 19743
rect 322 19641 356 19675
rect 322 19573 356 19607
rect 322 19505 356 19539
rect 322 19437 356 19471
rect 322 19369 356 19403
rect 322 19301 356 19335
rect 322 19233 356 19267
rect 322 19165 356 19199
rect 322 19097 356 19131
rect 322 19029 356 19063
rect 322 18961 356 18995
rect 322 18893 356 18927
rect 322 18825 356 18859
rect 322 18757 356 18791
rect 322 18689 356 18723
rect 322 18621 356 18655
rect 322 18553 356 18587
rect 322 18485 356 18519
rect 322 18417 356 18451
rect 322 18349 356 18383
rect 322 18281 356 18315
rect 322 18213 356 18247
rect 322 18145 356 18179
rect 322 18077 356 18111
rect 322 18009 356 18043
rect 322 17941 356 17975
rect 322 17873 356 17907
rect 322 17805 356 17839
rect 322 17737 356 17771
rect 322 17669 356 17703
rect 322 17601 356 17635
rect 322 17533 356 17567
rect 322 17465 356 17499
rect 322 17397 356 17431
rect 322 17329 356 17363
rect 322 17261 356 17295
rect 322 17193 356 17227
rect 322 17125 356 17159
rect 322 17057 356 17091
rect 322 16989 356 17023
rect 322 16921 356 16955
rect 322 16853 356 16887
rect 322 16785 356 16819
rect 322 16717 356 16751
rect 322 16649 356 16683
rect 322 16581 356 16615
rect 322 16513 356 16547
rect 322 16445 356 16479
rect 322 16377 356 16411
rect 322 16309 356 16343
rect 322 16241 356 16275
rect 322 16173 356 16207
rect 322 16105 356 16139
rect 322 16037 356 16071
rect 322 15969 356 16003
rect 322 15901 356 15935
rect 322 15833 356 15867
rect 322 15765 356 15799
rect 322 15697 356 15731
rect 322 15629 356 15663
rect 322 15561 356 15595
rect 322 15493 356 15527
rect 322 15425 356 15459
rect 322 15357 356 15391
rect 322 15289 356 15323
rect 322 15221 356 15255
rect 322 15153 356 15187
rect 322 15085 356 15119
rect 322 15017 356 15051
rect 322 14949 356 14983
rect 322 14881 356 14915
rect 322 14813 356 14847
rect 322 14745 356 14779
rect 322 14677 356 14711
rect 322 14609 356 14643
rect 322 14541 356 14575
rect 322 14473 356 14507
rect 322 14405 356 14439
rect 322 14337 356 14371
rect 322 14269 356 14303
rect 322 14201 356 14235
rect 322 14133 356 14167
rect 322 14065 356 14099
rect 322 13997 356 14031
rect 322 13929 356 13963
rect 322 13861 356 13895
rect 322 13793 356 13827
rect 322 13725 356 13759
rect 322 13657 356 13691
rect 322 13589 356 13623
rect 322 13521 356 13555
rect 322 13453 356 13487
rect 322 13385 356 13419
rect 322 13317 356 13351
rect 322 13249 356 13283
rect 322 13181 356 13215
rect 322 13113 356 13147
rect 322 13045 356 13079
rect 322 12977 356 13011
rect 322 12909 356 12943
rect 322 12841 356 12875
rect 322 12773 356 12807
rect 322 12705 356 12739
rect 322 12637 356 12671
rect 322 12569 356 12603
rect 322 12501 356 12535
rect 322 12433 356 12467
rect 322 12365 356 12399
rect 322 12297 356 12331
rect 322 12229 356 12263
rect 322 12161 356 12195
rect 322 12093 356 12127
rect 322 12025 356 12059
rect 322 11957 356 11991
rect 322 11889 356 11923
rect 322 11821 356 11855
rect 322 11753 356 11787
rect 322 11685 356 11719
rect 322 11617 356 11651
rect 322 11549 356 11583
rect 322 11481 356 11515
rect 322 11413 356 11447
rect 322 11345 356 11379
rect 322 11277 356 11311
rect 322 11209 356 11243
rect 322 11141 356 11175
rect 322 11073 356 11107
rect 322 11005 356 11039
rect 322 10937 356 10971
rect 322 10869 356 10903
rect 322 10801 356 10835
rect 322 10733 356 10767
rect 322 10665 356 10699
rect 322 10597 356 10631
rect 322 10529 356 10563
rect 322 10461 356 10495
rect 322 10393 356 10427
rect 322 10325 356 10359
rect 322 10257 356 10291
rect 322 10189 356 10223
rect 322 10121 356 10155
rect 322 10053 356 10087
rect 322 9985 356 10019
rect 322 9917 356 9951
rect 322 9849 356 9883
rect 322 9781 356 9815
rect 322 9713 356 9747
rect 1365 34602 1399 34636
rect 1433 34602 1467 34636
rect 1501 34602 1535 34636
rect 1569 34602 1603 34636
rect 1637 34602 1671 34636
rect 1705 34602 1739 34636
rect 1773 34602 1807 34636
rect 1841 34602 1875 34636
rect 1909 34602 1943 34636
rect 1977 34602 2011 34636
rect 2045 34602 2079 34636
rect 2113 34602 2147 34636
rect 2181 34602 2215 34636
rect 2249 34602 2283 34636
rect 2317 34602 2351 34636
rect 2385 34602 2419 34636
rect 2453 34602 2487 34636
rect 2521 34602 2555 34636
rect 2589 34602 2623 34636
rect 2657 34602 2691 34636
rect 2725 34602 2759 34636
rect 2793 34602 2827 34636
rect 2861 34602 2895 34636
rect 2929 34602 2963 34636
rect 2997 34602 3031 34636
rect 3065 34602 3099 34636
rect 3133 34602 3167 34636
rect 3201 34602 3235 34636
rect 3269 34602 3303 34636
rect 3337 34602 3371 34636
rect 3405 34602 3439 34636
rect 3473 34602 3507 34636
rect 3541 34602 3575 34636
rect 3609 34602 3643 34636
rect 3677 34602 3711 34636
rect 3745 34602 3779 34636
rect 3813 34602 3847 34636
rect 3881 34602 3915 34636
rect 3949 34602 3983 34636
rect 4017 34602 4051 34636
rect 4085 34602 4119 34636
rect 4153 34602 4187 34636
rect 4221 34602 4255 34636
rect 4289 34602 4323 34636
rect 4357 34602 4391 34636
rect 4425 34602 4459 34636
rect 4493 34602 4527 34636
rect 4561 34602 4595 34636
rect 4629 34602 4663 34636
rect 4697 34602 4731 34636
rect 4765 34602 4799 34636
rect 4833 34602 4867 34636
rect 4901 34602 4935 34636
rect 4969 34602 5003 34636
rect 5037 34602 5071 34636
rect 5105 34602 5139 34636
rect 5173 34602 5207 34636
rect 5241 34602 5275 34636
rect 5309 34602 5343 34636
rect 5377 34602 5411 34636
rect 5445 34602 5479 34636
rect 5513 34602 5547 34636
rect 5581 34602 5615 34636
rect 5649 34602 5683 34636
rect 5717 34602 5751 34636
rect 5785 34602 5819 34636
rect 5853 34602 5887 34636
rect 5921 34602 5955 34636
rect 5989 34602 6023 34636
rect 6057 34602 6091 34636
rect 6125 34602 6159 34636
rect 6193 34602 6227 34636
rect 6261 34602 6295 34636
rect 6329 34602 6363 34636
rect 6397 34602 6431 34636
rect 6465 34602 6499 34636
rect 6533 34602 6567 34636
rect 6601 34602 6635 34636
rect 6669 34602 6703 34636
rect 6737 34602 6771 34636
rect 6805 34602 6839 34636
rect 6873 34602 6907 34636
rect 6941 34602 6975 34636
rect 7009 34602 7043 34636
rect 7077 34602 7111 34636
rect 7145 34602 7179 34636
rect 7213 34602 7247 34636
rect 7281 34602 7315 34636
rect 7349 34602 7383 34636
rect 7417 34602 7451 34636
rect 7485 34602 7519 34636
rect 7553 34602 7587 34636
rect 7621 34602 7655 34636
rect 7689 34602 7723 34636
rect 7757 34602 7791 34636
rect 7825 34602 7859 34636
rect 7893 34602 7927 34636
rect 7961 34602 7995 34636
rect 8029 34602 8063 34636
rect 8097 34602 8131 34636
rect 8165 34602 8199 34636
rect 8233 34602 8267 34636
rect 8301 34602 8335 34636
rect 8369 34602 8403 34636
rect 8437 34602 8471 34636
rect 8505 34602 8539 34636
rect 8573 34602 8607 34636
rect 8641 34602 8675 34636
rect 8709 34602 8743 34636
rect 8777 34602 8811 34636
rect 8845 34602 8879 34636
rect 8913 34602 8947 34636
rect 8981 34602 9015 34636
rect 9049 34602 9083 34636
rect 9117 34602 9151 34636
rect 9185 34602 9219 34636
rect 9253 34602 9287 34636
rect 9321 34602 9355 34636
rect 9389 34602 9423 34636
rect 9457 34602 9491 34636
rect 9525 34602 9559 34636
rect 9593 34602 9627 34636
rect 9661 34602 9695 34636
rect 9729 34602 9763 34636
rect 9797 34602 9831 34636
rect 9865 34602 9899 34636
rect 9933 34602 9967 34636
rect 10001 34602 10035 34636
rect 10069 34602 10103 34636
rect 10137 34602 10171 34636
rect 10205 34602 10239 34636
rect 10273 34602 10307 34636
rect 10341 34602 10375 34636
rect 10409 34602 10443 34636
rect 10477 34602 10511 34636
rect 10545 34602 10579 34636
rect 10613 34602 10647 34636
rect 10681 34602 10715 34636
rect 10749 34602 10783 34636
rect 10817 34602 10851 34636
rect 10885 34602 10919 34636
rect 10953 34602 10987 34636
rect 11021 34602 11055 34636
rect 11089 34602 11123 34636
rect 11157 34602 11191 34636
rect 11225 34602 11259 34636
rect 11293 34602 11327 34636
rect 11361 34602 11395 34636
rect 11429 34602 11463 34636
rect 11497 34602 11531 34636
rect 11565 34602 11599 34636
rect 11633 34602 11667 34636
rect 11701 34602 11735 34636
rect 11769 34602 11803 34636
rect 11837 34602 11871 34636
rect 11905 34602 11939 34636
rect 11973 34602 12007 34636
rect 12041 34602 12075 34636
rect 12109 34602 12143 34636
rect 12177 34602 12211 34636
rect 12245 34602 12279 34636
rect 12313 34602 12347 34636
rect 12381 34602 12415 34636
rect 12449 34602 12483 34636
rect 12517 34602 12551 34636
rect 12585 34602 12619 34636
rect 12653 34602 12687 34636
rect 12721 34602 12755 34636
rect 12789 34602 12823 34636
rect 12857 34602 12891 34636
rect 12925 34602 12959 34636
rect 12993 34602 13027 34636
rect 13061 34602 13095 34636
rect 13129 34602 13163 34636
rect 13197 34602 13231 34636
rect 13265 34602 13299 34636
rect 13333 34602 13367 34636
rect 13401 34602 13435 34636
rect 13469 34602 13503 34636
rect 13537 34602 13571 34636
rect 13605 34602 13639 34636
rect 1221 34452 1255 34486
rect 1221 34384 1255 34418
rect 1221 34316 1255 34350
rect 1221 34248 1255 34282
rect 1221 34180 1255 34214
rect 1221 34112 1255 34146
rect 1221 34044 1255 34078
rect 1221 33976 1255 34010
rect 1221 33908 1255 33942
rect 1221 33840 1255 33874
rect 1221 33772 1255 33806
rect 1221 33704 1255 33738
rect 1221 33636 1255 33670
rect 1221 33568 1255 33602
rect 1221 33500 1255 33534
rect 1221 33432 1255 33466
rect 1221 33364 1255 33398
rect 1221 33296 1255 33330
rect 1221 33228 1255 33262
rect 1221 33160 1255 33194
rect 1221 33092 1255 33126
rect 1221 33024 1255 33058
rect 1221 32956 1255 32990
rect 1221 32888 1255 32922
rect 1221 32820 1255 32854
rect 1221 32752 1255 32786
rect 1221 32684 1255 32718
rect 1221 32616 1255 32650
rect 1221 32548 1255 32582
rect 1221 32480 1255 32514
rect 1221 32412 1255 32446
rect 1221 32344 1255 32378
rect 1221 32276 1255 32310
rect 1221 32208 1255 32242
rect 1221 32140 1255 32174
rect 1221 32072 1255 32106
rect 1221 32004 1255 32038
rect 1221 31936 1255 31970
rect 1221 31868 1255 31902
rect 1221 31800 1255 31834
rect 1221 31732 1255 31766
rect 1221 31664 1255 31698
rect 1221 31596 1255 31630
rect 1221 31528 1255 31562
rect 1221 31460 1255 31494
rect 1221 31392 1255 31426
rect 1221 31324 1255 31358
rect 1221 31256 1255 31290
rect 1221 31188 1255 31222
rect 1221 31120 1255 31154
rect 1221 31052 1255 31086
rect 1221 30984 1255 31018
rect 1221 30916 1255 30950
rect 1221 30848 1255 30882
rect 1221 30780 1255 30814
rect 1221 30712 1255 30746
rect 1221 30644 1255 30678
rect 1221 30576 1255 30610
rect 1221 30508 1255 30542
rect 1221 30440 1255 30474
rect 1221 30372 1255 30406
rect 1221 30304 1255 30338
rect 1221 30236 1255 30270
rect 1221 30168 1255 30202
rect 1221 30100 1255 30134
rect 1221 30032 1255 30066
rect 1221 29964 1255 29998
rect 1221 29896 1255 29930
rect 1221 29828 1255 29862
rect 1221 29760 1255 29794
rect 1221 29692 1255 29726
rect 1221 29624 1255 29658
rect 1221 29556 1255 29590
rect 1221 29488 1255 29522
rect 1221 29420 1255 29454
rect 1221 29352 1255 29386
rect 1221 29284 1255 29318
rect 1221 29216 1255 29250
rect 1221 29148 1255 29182
rect 1221 29080 1255 29114
rect 1221 29012 1255 29046
rect 1221 28944 1255 28978
rect 1221 28876 1255 28910
rect 1221 28808 1255 28842
rect 1221 28740 1255 28774
rect 1221 28672 1255 28706
rect 1221 28604 1255 28638
rect 1221 28536 1255 28570
rect 1221 28468 1255 28502
rect 1221 28400 1255 28434
rect 1221 28332 1255 28366
rect 1221 28264 1255 28298
rect 1221 28196 1255 28230
rect 1221 28128 1255 28162
rect 1221 28060 1255 28094
rect 1221 27992 1255 28026
rect 1221 27924 1255 27958
rect 1221 27856 1255 27890
rect 1221 27788 1255 27822
rect 1221 27720 1255 27754
rect 1221 27652 1255 27686
rect 1221 27584 1255 27618
rect 1221 27516 1255 27550
rect 1221 27448 1255 27482
rect 1221 27380 1255 27414
rect 1221 27312 1255 27346
rect 1221 27244 1255 27278
rect 1221 27176 1255 27210
rect 1221 27108 1255 27142
rect 1221 27040 1255 27074
rect 1221 26972 1255 27006
rect 1221 26904 1255 26938
rect 1221 26836 1255 26870
rect 1221 26768 1255 26802
rect 1221 26700 1255 26734
rect 1221 26632 1255 26666
rect 1221 26564 1255 26598
rect 1221 26496 1255 26530
rect 1221 26428 1255 26462
rect 1221 26360 1255 26394
rect 1221 26292 1255 26326
rect 1221 26224 1255 26258
rect 1221 26156 1255 26190
rect 1221 26088 1255 26122
rect 1221 26020 1255 26054
rect 1221 25952 1255 25986
rect 1221 25884 1255 25918
rect 1221 25816 1255 25850
rect 1221 25748 1255 25782
rect 1221 25680 1255 25714
rect 1221 25612 1255 25646
rect 1221 25544 1255 25578
rect 1221 25476 1255 25510
rect 1221 25408 1255 25442
rect 1221 25340 1255 25374
rect 1221 25272 1255 25306
rect 1221 25204 1255 25238
rect 1221 25136 1255 25170
rect 1221 25068 1255 25102
rect 1221 25000 1255 25034
rect 1221 24932 1255 24966
rect 1221 24864 1255 24898
rect 1221 24796 1255 24830
rect 1221 24728 1255 24762
rect 1221 24660 1255 24694
rect 1221 24592 1255 24626
rect 1221 24524 1255 24558
rect 1221 24456 1255 24490
rect 1221 24388 1255 24422
rect 1221 24320 1255 24354
rect 1221 24252 1255 24286
rect 1221 24184 1255 24218
rect 1221 24116 1255 24150
rect 1221 24048 1255 24082
rect 1221 23980 1255 24014
rect 1221 23912 1255 23946
rect 1221 23844 1255 23878
rect 1221 23776 1255 23810
rect 1221 23708 1255 23742
rect 1221 23640 1255 23674
rect 1221 23572 1255 23606
rect 1221 23504 1255 23538
rect 1221 23436 1255 23470
rect 1221 23368 1255 23402
rect 1221 23300 1255 23334
rect 1221 23232 1255 23266
rect 1221 23164 1255 23198
rect 1221 23096 1255 23130
rect 1221 23028 1255 23062
rect 1221 22960 1255 22994
rect 1221 22892 1255 22926
rect 1221 22824 1255 22858
rect 1221 22756 1255 22790
rect 1221 22688 1255 22722
rect 1221 22620 1255 22654
rect 1221 22552 1255 22586
rect 1221 22484 1255 22518
rect 1221 22416 1255 22450
rect 1221 22348 1255 22382
rect 1221 22280 1255 22314
rect 1221 22212 1255 22246
rect 1221 22144 1255 22178
rect 1221 22076 1255 22110
rect 1221 22008 1255 22042
rect 1221 21940 1255 21974
rect 1221 21872 1255 21906
rect 1221 21804 1255 21838
rect 1221 21736 1255 21770
rect 1221 21668 1255 21702
rect 1221 21600 1255 21634
rect 1221 21532 1255 21566
rect 1221 21464 1255 21498
rect 1221 21396 1255 21430
rect 1221 21328 1255 21362
rect 1221 21260 1255 21294
rect 1221 21192 1255 21226
rect 1221 21124 1255 21158
rect 1221 21056 1255 21090
rect 1221 20988 1255 21022
rect 1221 20920 1255 20954
rect 1221 20852 1255 20886
rect 1221 20784 1255 20818
rect 1221 20716 1255 20750
rect 1221 20648 1255 20682
rect 1221 20580 1255 20614
rect 1221 20512 1255 20546
rect 1221 20444 1255 20478
rect 1221 20376 1255 20410
rect 1221 20308 1255 20342
rect 1221 20240 1255 20274
rect 1221 20172 1255 20206
rect 1221 20104 1255 20138
rect 1221 20036 1255 20070
rect 1221 19968 1255 20002
rect 1221 19900 1255 19934
rect 1221 19832 1255 19866
rect 1221 19764 1255 19798
rect 1221 19696 1255 19730
rect 1221 19628 1255 19662
rect 1221 19560 1255 19594
rect 1221 19492 1255 19526
rect 1221 19424 1255 19458
rect 1221 19356 1255 19390
rect 1221 19288 1255 19322
rect 1221 19220 1255 19254
rect 1221 19152 1255 19186
rect 1221 19084 1255 19118
rect 1221 19016 1255 19050
rect 1221 18948 1255 18982
rect 1221 18880 1255 18914
rect 1221 18812 1255 18846
rect 1221 18744 1255 18778
rect 1221 18676 1255 18710
rect 1221 18608 1255 18642
rect 1221 18540 1255 18574
rect 1221 18472 1255 18506
rect 1221 18404 1255 18438
rect 1221 18336 1255 18370
rect 1221 18268 1255 18302
rect 1221 18200 1255 18234
rect 1221 18132 1255 18166
rect 1221 18064 1255 18098
rect 1221 17996 1255 18030
rect 1221 17928 1255 17962
rect 1221 17860 1255 17894
rect 1221 17792 1255 17826
rect 1221 17724 1255 17758
rect 1221 17656 1255 17690
rect 1221 17588 1255 17622
rect 1221 17520 1255 17554
rect 1221 17452 1255 17486
rect 1221 17384 1255 17418
rect 1221 17316 1255 17350
rect 1221 17248 1255 17282
rect 1221 17180 1255 17214
rect 1221 17112 1255 17146
rect 1221 17044 1255 17078
rect 1221 16976 1255 17010
rect 1221 16908 1255 16942
rect 1221 16840 1255 16874
rect 1221 16772 1255 16806
rect 1221 16704 1255 16738
rect 1221 16636 1255 16670
rect 1221 16568 1255 16602
rect 1221 16500 1255 16534
rect 1221 16432 1255 16466
rect 1221 16364 1255 16398
rect 1221 16296 1255 16330
rect 1221 16228 1255 16262
rect 1221 16160 1255 16194
rect 1221 16092 1255 16126
rect 1221 16024 1255 16058
rect 1221 15956 1255 15990
rect 1221 15888 1255 15922
rect 1221 15820 1255 15854
rect 1221 15752 1255 15786
rect 1221 15684 1255 15718
rect 1221 15616 1255 15650
rect 1221 15548 1255 15582
rect 1221 15480 1255 15514
rect 1221 15412 1255 15446
rect 1221 15344 1255 15378
rect 1221 15276 1255 15310
rect 1221 15208 1255 15242
rect 1221 15140 1255 15174
rect 1221 15072 1255 15106
rect 1221 15004 1255 15038
rect 1221 14936 1255 14970
rect 1221 14868 1255 14902
rect 1221 14800 1255 14834
rect 1221 14732 1255 14766
rect 1221 14664 1255 14698
rect 1221 14596 1255 14630
rect 1221 14528 1255 14562
rect 1221 14460 1255 14494
rect 1221 14392 1255 14426
rect 1221 14324 1255 14358
rect 1221 14256 1255 14290
rect 1221 14188 1255 14222
rect 1221 14120 1255 14154
rect 1221 14052 1255 14086
rect 1221 13984 1255 14018
rect 1221 13916 1255 13950
rect 1221 13848 1255 13882
rect 1221 13780 1255 13814
rect 1221 13712 1255 13746
rect 1221 13644 1255 13678
rect 1221 13576 1255 13610
rect 1221 13508 1255 13542
rect 1221 13440 1255 13474
rect 1221 13372 1255 13406
rect 1221 13304 1255 13338
rect 1221 13236 1255 13270
rect 1221 13168 1255 13202
rect 1221 13100 1255 13134
rect 1221 13032 1255 13066
rect 1221 12964 1255 12998
rect 1221 12896 1255 12930
rect 1221 12828 1255 12862
rect 1221 12760 1255 12794
rect 1221 12692 1255 12726
rect 1221 12624 1255 12658
rect 1221 12556 1255 12590
rect 1221 12488 1255 12522
rect 1221 12420 1255 12454
rect 1221 12352 1255 12386
rect 1221 12284 1255 12318
rect 1221 12216 1255 12250
rect 1221 12148 1255 12182
rect 1221 12080 1255 12114
rect 1221 12012 1255 12046
rect 1221 11944 1255 11978
rect 1221 11876 1255 11910
rect 1221 11808 1255 11842
rect 1221 11740 1255 11774
rect 1221 11672 1255 11706
rect 1221 11604 1255 11638
rect 1221 11536 1255 11570
rect 1221 11468 1255 11502
rect 1221 11400 1255 11434
rect 1221 11332 1255 11366
rect 1221 11264 1255 11298
rect 1221 11196 1255 11230
rect 1221 11128 1255 11162
rect 1221 11060 1255 11094
rect 1221 10992 1255 11026
rect 1221 10924 1255 10958
rect 1221 10856 1255 10890
rect 1221 10788 1255 10822
rect 1221 10720 1255 10754
rect 1221 10652 1255 10686
rect 1221 10584 1255 10618
rect 1221 10516 1255 10550
rect 1221 10448 1255 10482
rect 1221 10380 1255 10414
rect 13739 34456 13773 34490
rect 13739 34388 13773 34422
rect 13739 34320 13773 34354
rect 13739 34252 13773 34286
rect 13739 34184 13773 34218
rect 13739 34116 13773 34150
rect 13739 34048 13773 34082
rect 13739 33980 13773 34014
rect 13739 33912 13773 33946
rect 13739 33844 13773 33878
rect 13739 33776 13773 33810
rect 13739 33708 13773 33742
rect 13739 33640 13773 33674
rect 13739 33572 13773 33606
rect 13739 33504 13773 33538
rect 13739 33436 13773 33470
rect 13739 33368 13773 33402
rect 13739 33300 13773 33334
rect 13739 33232 13773 33266
rect 13739 33164 13773 33198
rect 13739 33096 13773 33130
rect 13739 33028 13773 33062
rect 13739 32960 13773 32994
rect 13739 32892 13773 32926
rect 13739 32824 13773 32858
rect 13739 32756 13773 32790
rect 13739 32688 13773 32722
rect 13739 32620 13773 32654
rect 13739 32552 13773 32586
rect 13739 32484 13773 32518
rect 13739 32416 13773 32450
rect 13739 32348 13773 32382
rect 13739 32280 13773 32314
rect 13739 32212 13773 32246
rect 13739 32144 13773 32178
rect 13739 32076 13773 32110
rect 13739 32008 13773 32042
rect 13739 31940 13773 31974
rect 13739 31872 13773 31906
rect 13739 31804 13773 31838
rect 13739 31736 13773 31770
rect 13739 31668 13773 31702
rect 13739 31600 13773 31634
rect 13739 31532 13773 31566
rect 13739 31464 13773 31498
rect 13739 31396 13773 31430
rect 13739 31328 13773 31362
rect 13739 31260 13773 31294
rect 13739 31192 13773 31226
rect 13739 31124 13773 31158
rect 13739 31056 13773 31090
rect 13739 30988 13773 31022
rect 13739 30920 13773 30954
rect 13739 30852 13773 30886
rect 13739 30784 13773 30818
rect 13739 30716 13773 30750
rect 13739 30648 13773 30682
rect 13739 30580 13773 30614
rect 13739 30512 13773 30546
rect 13739 30444 13773 30478
rect 13739 30376 13773 30410
rect 13739 30308 13773 30342
rect 13739 30240 13773 30274
rect 13739 30172 13773 30206
rect 13739 30104 13773 30138
rect 13739 30036 13773 30070
rect 13739 29968 13773 30002
rect 13739 29900 13773 29934
rect 13739 29832 13773 29866
rect 13739 29764 13773 29798
rect 13739 29696 13773 29730
rect 13739 29628 13773 29662
rect 13739 29560 13773 29594
rect 13739 29492 13773 29526
rect 13739 29424 13773 29458
rect 13739 29356 13773 29390
rect 13739 29288 13773 29322
rect 13739 29220 13773 29254
rect 13739 29152 13773 29186
rect 13739 29084 13773 29118
rect 13739 29016 13773 29050
rect 13739 28948 13773 28982
rect 13739 28880 13773 28914
rect 13739 28812 13773 28846
rect 13739 28744 13773 28778
rect 13739 28676 13773 28710
rect 13739 28608 13773 28642
rect 13739 28540 13773 28574
rect 13739 28472 13773 28506
rect 13739 28404 13773 28438
rect 13739 28336 13773 28370
rect 13739 28268 13773 28302
rect 13739 28200 13773 28234
rect 13739 28132 13773 28166
rect 13739 28064 13773 28098
rect 13739 27996 13773 28030
rect 13739 27928 13773 27962
rect 13739 27860 13773 27894
rect 13739 27792 13773 27826
rect 13739 27724 13773 27758
rect 13739 27656 13773 27690
rect 13739 27588 13773 27622
rect 13739 27520 13773 27554
rect 13739 27452 13773 27486
rect 13739 27384 13773 27418
rect 13739 27316 13773 27350
rect 13739 27248 13773 27282
rect 13739 27180 13773 27214
rect 13739 27112 13773 27146
rect 13739 27044 13773 27078
rect 13739 26976 13773 27010
rect 13739 26908 13773 26942
rect 13739 26840 13773 26874
rect 13739 26772 13773 26806
rect 13739 26704 13773 26738
rect 13739 26636 13773 26670
rect 13739 26568 13773 26602
rect 13739 26500 13773 26534
rect 13739 26432 13773 26466
rect 13739 26364 13773 26398
rect 13739 26296 13773 26330
rect 13739 26228 13773 26262
rect 13739 26160 13773 26194
rect 13739 26092 13773 26126
rect 13739 26024 13773 26058
rect 13739 25956 13773 25990
rect 13739 25888 13773 25922
rect 13739 25820 13773 25854
rect 13739 25752 13773 25786
rect 13739 25684 13773 25718
rect 13739 25616 13773 25650
rect 13739 25548 13773 25582
rect 13739 25480 13773 25514
rect 13739 25412 13773 25446
rect 13739 25344 13773 25378
rect 13739 25276 13773 25310
rect 13739 25208 13773 25242
rect 13739 25140 13773 25174
rect 13739 25072 13773 25106
rect 13739 25004 13773 25038
rect 13739 24936 13773 24970
rect 13739 24868 13773 24902
rect 13739 24800 13773 24834
rect 13739 24732 13773 24766
rect 13739 24664 13773 24698
rect 13739 24596 13773 24630
rect 13739 24528 13773 24562
rect 13739 24460 13773 24494
rect 13739 24392 13773 24426
rect 13739 24324 13773 24358
rect 13739 24256 13773 24290
rect 13739 24188 13773 24222
rect 13739 24120 13773 24154
rect 13739 24052 13773 24086
rect 13739 23984 13773 24018
rect 13739 23916 13773 23950
rect 13739 23848 13773 23882
rect 13739 23780 13773 23814
rect 13739 23712 13773 23746
rect 13739 23644 13773 23678
rect 13739 23576 13773 23610
rect 13739 23508 13773 23542
rect 13739 23440 13773 23474
rect 13739 23372 13773 23406
rect 13739 23304 13773 23338
rect 13739 23236 13773 23270
rect 13739 23168 13773 23202
rect 13739 23100 13773 23134
rect 13739 23032 13773 23066
rect 13739 22964 13773 22998
rect 13739 22896 13773 22930
rect 13739 22828 13773 22862
rect 13739 22760 13773 22794
rect 13739 22692 13773 22726
rect 13739 22624 13773 22658
rect 13739 22556 13773 22590
rect 13739 22488 13773 22522
rect 13739 22420 13773 22454
rect 13739 22352 13773 22386
rect 13739 22284 13773 22318
rect 13739 22216 13773 22250
rect 13739 22148 13773 22182
rect 13739 22080 13773 22114
rect 13739 22012 13773 22046
rect 13739 21944 13773 21978
rect 13739 21876 13773 21910
rect 13739 21808 13773 21842
rect 13739 21740 13773 21774
rect 13739 21672 13773 21706
rect 13739 21604 13773 21638
rect 13739 21536 13773 21570
rect 13739 21468 13773 21502
rect 13739 21400 13773 21434
rect 13739 21332 13773 21366
rect 13739 21264 13773 21298
rect 13739 21196 13773 21230
rect 13739 21128 13773 21162
rect 13739 21060 13773 21094
rect 13739 20992 13773 21026
rect 13739 20924 13773 20958
rect 13739 20856 13773 20890
rect 13739 20788 13773 20822
rect 13739 20720 13773 20754
rect 13739 20652 13773 20686
rect 13739 20584 13773 20618
rect 13739 20516 13773 20550
rect 13739 20448 13773 20482
rect 13739 20380 13773 20414
rect 13739 20312 13773 20346
rect 13739 20244 13773 20278
rect 13739 20176 13773 20210
rect 13739 20108 13773 20142
rect 13739 20040 13773 20074
rect 13739 19972 13773 20006
rect 13739 19904 13773 19938
rect 13739 19836 13773 19870
rect 13739 19768 13773 19802
rect 13739 19700 13773 19734
rect 13739 19632 13773 19666
rect 13739 19564 13773 19598
rect 13739 19496 13773 19530
rect 13739 19428 13773 19462
rect 13739 19360 13773 19394
rect 13739 19292 13773 19326
rect 13739 19224 13773 19258
rect 13739 19156 13773 19190
rect 13739 19088 13773 19122
rect 13739 19020 13773 19054
rect 13739 18952 13773 18986
rect 13739 18884 13773 18918
rect 13739 18816 13773 18850
rect 13739 18748 13773 18782
rect 13739 18680 13773 18714
rect 13739 18612 13773 18646
rect 13739 18544 13773 18578
rect 13739 18476 13773 18510
rect 13739 18408 13773 18442
rect 13739 18340 13773 18374
rect 13739 18272 13773 18306
rect 13739 18204 13773 18238
rect 13739 18136 13773 18170
rect 13739 18068 13773 18102
rect 13739 18000 13773 18034
rect 13739 17932 13773 17966
rect 13739 17864 13773 17898
rect 13739 17796 13773 17830
rect 13739 17728 13773 17762
rect 13739 17660 13773 17694
rect 13739 17592 13773 17626
rect 13739 17524 13773 17558
rect 13739 17456 13773 17490
rect 13739 17388 13773 17422
rect 13739 17320 13773 17354
rect 13739 17252 13773 17286
rect 13739 17184 13773 17218
rect 13739 17116 13773 17150
rect 13739 17048 13773 17082
rect 13739 16980 13773 17014
rect 13739 16912 13773 16946
rect 13739 16844 13773 16878
rect 13739 16776 13773 16810
rect 13739 16708 13773 16742
rect 13739 16640 13773 16674
rect 13739 16572 13773 16606
rect 13739 16504 13773 16538
rect 13739 16436 13773 16470
rect 13739 16368 13773 16402
rect 13739 16300 13773 16334
rect 13739 16232 13773 16266
rect 13739 16164 13773 16198
rect 13739 16096 13773 16130
rect 13739 16028 13773 16062
rect 13739 15960 13773 15994
rect 13739 15892 13773 15926
rect 13739 15824 13773 15858
rect 13739 15756 13773 15790
rect 13739 15688 13773 15722
rect 13739 15620 13773 15654
rect 13739 15552 13773 15586
rect 13739 15484 13773 15518
rect 13739 15416 13773 15450
rect 13739 15348 13773 15382
rect 13739 15280 13773 15314
rect 13739 15212 13773 15246
rect 13739 15144 13773 15178
rect 13739 15076 13773 15110
rect 13739 15008 13773 15042
rect 13739 14940 13773 14974
rect 13739 14872 13773 14906
rect 13739 14804 13773 14838
rect 13739 14736 13773 14770
rect 13739 14668 13773 14702
rect 13739 14600 13773 14634
rect 13739 14532 13773 14566
rect 13739 14464 13773 14498
rect 13739 14396 13773 14430
rect 13739 14328 13773 14362
rect 13739 14260 13773 14294
rect 13739 14192 13773 14226
rect 13739 14124 13773 14158
rect 13739 14056 13773 14090
rect 13739 13988 13773 14022
rect 13739 13920 13773 13954
rect 13739 13852 13773 13886
rect 13739 13784 13773 13818
rect 13739 13716 13773 13750
rect 13739 13648 13773 13682
rect 13739 13580 13773 13614
rect 13739 13512 13773 13546
rect 13739 13444 13773 13478
rect 13739 13376 13773 13410
rect 13739 13308 13773 13342
rect 13739 13240 13773 13274
rect 13739 13172 13773 13206
rect 13739 13104 13773 13138
rect 13739 13036 13773 13070
rect 13739 12968 13773 13002
rect 13739 12900 13773 12934
rect 13739 12832 13773 12866
rect 13739 12764 13773 12798
rect 13739 12696 13773 12730
rect 13739 12628 13773 12662
rect 13739 12560 13773 12594
rect 13739 12492 13773 12526
rect 13739 12424 13773 12458
rect 13739 12356 13773 12390
rect 13739 12288 13773 12322
rect 13739 12220 13773 12254
rect 13739 12152 13773 12186
rect 13739 12084 13773 12118
rect 13739 12016 13773 12050
rect 13739 11948 13773 11982
rect 13739 11880 13773 11914
rect 13739 11812 13773 11846
rect 13739 11744 13773 11778
rect 13739 11676 13773 11710
rect 13739 11608 13773 11642
rect 13739 11540 13773 11574
rect 13739 11472 13773 11506
rect 13739 11404 13773 11438
rect 13739 11336 13773 11370
rect 13739 11268 13773 11302
rect 13739 11200 13773 11234
rect 13739 11132 13773 11166
rect 13739 11064 13773 11098
rect 13739 10996 13773 11030
rect 13739 10928 13773 10962
rect 13739 10860 13773 10894
rect 13739 10792 13773 10826
rect 13739 10724 13773 10758
rect 13739 10656 13773 10690
rect 13739 10588 13773 10622
rect 13739 10520 13773 10554
rect 13739 10452 13773 10486
rect 13739 10384 13773 10418
rect 1355 10256 1389 10290
rect 1423 10256 1457 10290
rect 1491 10256 1525 10290
rect 1559 10256 1593 10290
rect 1627 10256 1661 10290
rect 1695 10256 1729 10290
rect 1763 10256 1797 10290
rect 1831 10256 1865 10290
rect 1899 10256 1933 10290
rect 1967 10256 2001 10290
rect 2035 10256 2069 10290
rect 2103 10256 2137 10290
rect 2171 10256 2205 10290
rect 2239 10256 2273 10290
rect 2307 10256 2341 10290
rect 2375 10256 2409 10290
rect 2443 10256 2477 10290
rect 2511 10256 2545 10290
rect 2579 10256 2613 10290
rect 2647 10256 2681 10290
rect 2715 10256 2749 10290
rect 2783 10256 2817 10290
rect 2851 10256 2885 10290
rect 2919 10256 2953 10290
rect 2987 10256 3021 10290
rect 3055 10256 3089 10290
rect 3123 10256 3157 10290
rect 3191 10256 3225 10290
rect 3259 10256 3293 10290
rect 3327 10256 3361 10290
rect 3395 10256 3429 10290
rect 3463 10256 3497 10290
rect 3531 10256 3565 10290
rect 3599 10256 3633 10290
rect 3667 10256 3701 10290
rect 3735 10256 3769 10290
rect 3803 10256 3837 10290
rect 3871 10256 3905 10290
rect 3939 10256 3973 10290
rect 4007 10256 4041 10290
rect 4075 10256 4109 10290
rect 4143 10256 4177 10290
rect 4211 10256 4245 10290
rect 4279 10256 4313 10290
rect 4347 10256 4381 10290
rect 4415 10256 4449 10290
rect 4483 10256 4517 10290
rect 4551 10256 4585 10290
rect 4619 10256 4653 10290
rect 4687 10256 4721 10290
rect 4755 10256 4789 10290
rect 4823 10256 4857 10290
rect 4891 10256 4925 10290
rect 4959 10256 4993 10290
rect 5027 10256 5061 10290
rect 5095 10256 5129 10290
rect 5163 10256 5197 10290
rect 5231 10256 5265 10290
rect 5299 10256 5333 10290
rect 5367 10256 5401 10290
rect 5435 10256 5469 10290
rect 5503 10256 5537 10290
rect 5571 10256 5605 10290
rect 5639 10256 5673 10290
rect 5707 10256 5741 10290
rect 5775 10256 5809 10290
rect 5843 10256 5877 10290
rect 5911 10256 5945 10290
rect 5979 10256 6013 10290
rect 6047 10256 6081 10290
rect 6115 10256 6149 10290
rect 6183 10256 6217 10290
rect 6251 10256 6285 10290
rect 6319 10256 6353 10290
rect 6387 10256 6421 10290
rect 6455 10256 6489 10290
rect 6523 10256 6557 10290
rect 6591 10256 6625 10290
rect 6659 10256 6693 10290
rect 6727 10256 6761 10290
rect 6795 10256 6829 10290
rect 6863 10256 6897 10290
rect 6931 10256 6965 10290
rect 6999 10256 7033 10290
rect 7067 10256 7101 10290
rect 7135 10256 7169 10290
rect 7203 10256 7237 10290
rect 7271 10256 7305 10290
rect 7339 10256 7373 10290
rect 7407 10256 7441 10290
rect 7475 10256 7509 10290
rect 7543 10256 7577 10290
rect 7611 10256 7645 10290
rect 7679 10256 7713 10290
rect 7747 10256 7781 10290
rect 7815 10256 7849 10290
rect 7883 10256 7917 10290
rect 7951 10256 7985 10290
rect 8019 10256 8053 10290
rect 8087 10256 8121 10290
rect 8155 10256 8189 10290
rect 8223 10256 8257 10290
rect 8291 10256 8325 10290
rect 8359 10256 8393 10290
rect 8427 10256 8461 10290
rect 8495 10256 8529 10290
rect 8563 10256 8597 10290
rect 8631 10256 8665 10290
rect 8699 10256 8733 10290
rect 8767 10256 8801 10290
rect 8835 10256 8869 10290
rect 8903 10256 8937 10290
rect 8971 10256 9005 10290
rect 9039 10256 9073 10290
rect 9107 10256 9141 10290
rect 9175 10256 9209 10290
rect 9243 10256 9277 10290
rect 9311 10256 9345 10290
rect 9379 10256 9413 10290
rect 9447 10256 9481 10290
rect 9515 10256 9549 10290
rect 9583 10256 9617 10290
rect 9651 10256 9685 10290
rect 9719 10256 9753 10290
rect 9787 10256 9821 10290
rect 9855 10256 9889 10290
rect 9923 10256 9957 10290
rect 9991 10256 10025 10290
rect 10059 10256 10093 10290
rect 10127 10256 10161 10290
rect 10195 10256 10229 10290
rect 10263 10256 10297 10290
rect 10331 10256 10365 10290
rect 10399 10256 10433 10290
rect 10467 10256 10501 10290
rect 10535 10256 10569 10290
rect 10603 10256 10637 10290
rect 10671 10256 10705 10290
rect 10739 10256 10773 10290
rect 10807 10256 10841 10290
rect 10875 10256 10909 10290
rect 10943 10256 10977 10290
rect 11011 10256 11045 10290
rect 11079 10256 11113 10290
rect 11147 10256 11181 10290
rect 11215 10256 11249 10290
rect 11283 10256 11317 10290
rect 11351 10256 11385 10290
rect 11419 10256 11453 10290
rect 11487 10256 11521 10290
rect 11555 10256 11589 10290
rect 11623 10256 11657 10290
rect 11691 10256 11725 10290
rect 11759 10256 11793 10290
rect 11827 10256 11861 10290
rect 11895 10256 11929 10290
rect 11963 10256 11997 10290
rect 12031 10256 12065 10290
rect 12099 10256 12133 10290
rect 12167 10256 12201 10290
rect 12235 10256 12269 10290
rect 12303 10256 12337 10290
rect 12371 10256 12405 10290
rect 12439 10256 12473 10290
rect 12507 10256 12541 10290
rect 12575 10256 12609 10290
rect 12643 10256 12677 10290
rect 12711 10256 12745 10290
rect 12779 10256 12813 10290
rect 12847 10256 12881 10290
rect 12915 10256 12949 10290
rect 12983 10256 13017 10290
rect 13051 10256 13085 10290
rect 13119 10256 13153 10290
rect 13187 10256 13221 10290
rect 13255 10256 13289 10290
rect 13323 10256 13357 10290
rect 13391 10256 13425 10290
rect 13459 10256 13493 10290
rect 13527 10256 13561 10290
rect 13595 10256 13629 10290
rect 14609 36225 14643 36259
rect 14609 36157 14643 36191
rect 14609 36089 14643 36123
rect 14609 36021 14643 36055
rect 14609 35953 14643 35987
rect 14609 35885 14643 35919
rect 14609 35817 14643 35851
rect 14609 35749 14643 35783
rect 14609 35681 14643 35715
rect 14609 35613 14643 35647
rect 14609 35545 14643 35579
rect 14609 35477 14643 35511
rect 14609 35409 14643 35443
rect 14609 35341 14643 35375
rect 14609 35273 14643 35307
rect 14609 35205 14643 35239
rect 14609 35137 14643 35171
rect 14609 35069 14643 35103
rect 14609 35001 14643 35035
rect 14609 34933 14643 34967
rect 14609 34865 14643 34899
rect 14609 34797 14643 34831
rect 14609 34729 14643 34763
rect 14609 34661 14643 34695
rect 14609 34593 14643 34627
rect 14609 34525 14643 34559
rect 14609 34457 14643 34491
rect 14609 34389 14643 34423
rect 14609 34321 14643 34355
rect 14609 34253 14643 34287
rect 14609 34185 14643 34219
rect 14609 34117 14643 34151
rect 14609 34049 14643 34083
rect 14609 33981 14643 34015
rect 14609 33913 14643 33947
rect 14609 33845 14643 33879
rect 14609 33777 14643 33811
rect 14609 33709 14643 33743
rect 14609 33641 14643 33675
rect 14609 33573 14643 33607
rect 14609 33505 14643 33539
rect 14609 33437 14643 33471
rect 14609 33369 14643 33403
rect 14609 33301 14643 33335
rect 14609 33233 14643 33267
rect 14609 33165 14643 33199
rect 14609 33097 14643 33131
rect 14609 33029 14643 33063
rect 14609 32961 14643 32995
rect 14609 32893 14643 32927
rect 14609 32825 14643 32859
rect 14609 32757 14643 32791
rect 14609 32689 14643 32723
rect 14609 32621 14643 32655
rect 14609 32553 14643 32587
rect 14609 32485 14643 32519
rect 14609 32417 14643 32451
rect 14609 32349 14643 32383
rect 14609 32281 14643 32315
rect 14609 32213 14643 32247
rect 14609 32145 14643 32179
rect 14609 32077 14643 32111
rect 14609 32009 14643 32043
rect 14609 31941 14643 31975
rect 14609 31873 14643 31907
rect 14609 31805 14643 31839
rect 14609 31737 14643 31771
rect 14609 31669 14643 31703
rect 14609 31601 14643 31635
rect 14609 31533 14643 31567
rect 14609 31465 14643 31499
rect 14609 31397 14643 31431
rect 14609 31329 14643 31363
rect 14609 31261 14643 31295
rect 14609 31193 14643 31227
rect 14609 31125 14643 31159
rect 14609 31057 14643 31091
rect 14609 30989 14643 31023
rect 14609 30921 14643 30955
rect 14609 30853 14643 30887
rect 14609 30785 14643 30819
rect 14609 30717 14643 30751
rect 14609 30649 14643 30683
rect 14609 30581 14643 30615
rect 14609 30513 14643 30547
rect 14609 30445 14643 30479
rect 14609 30377 14643 30411
rect 14609 30309 14643 30343
rect 14609 30241 14643 30275
rect 14609 30173 14643 30207
rect 14609 30105 14643 30139
rect 14609 30037 14643 30071
rect 14609 29969 14643 30003
rect 14609 29901 14643 29935
rect 14609 29833 14643 29867
rect 14609 29765 14643 29799
rect 14609 29697 14643 29731
rect 14609 29629 14643 29663
rect 14609 29561 14643 29595
rect 14609 29493 14643 29527
rect 14609 29425 14643 29459
rect 14609 29357 14643 29391
rect 14609 29289 14643 29323
rect 14609 29221 14643 29255
rect 14609 29153 14643 29187
rect 14609 29085 14643 29119
rect 14609 29017 14643 29051
rect 14609 28949 14643 28983
rect 14609 28881 14643 28915
rect 14609 28813 14643 28847
rect 14609 28745 14643 28779
rect 14609 28677 14643 28711
rect 14609 28609 14643 28643
rect 14609 28541 14643 28575
rect 14609 28473 14643 28507
rect 14609 28405 14643 28439
rect 14609 28337 14643 28371
rect 14609 28269 14643 28303
rect 14609 28201 14643 28235
rect 14609 28133 14643 28167
rect 14609 28065 14643 28099
rect 14609 27997 14643 28031
rect 14609 27929 14643 27963
rect 14609 27861 14643 27895
rect 14609 27793 14643 27827
rect 14609 27725 14643 27759
rect 14609 27657 14643 27691
rect 14609 27589 14643 27623
rect 14609 27521 14643 27555
rect 14609 27453 14643 27487
rect 14609 27385 14643 27419
rect 14609 27317 14643 27351
rect 14609 27249 14643 27283
rect 14609 27181 14643 27215
rect 14609 27113 14643 27147
rect 14609 27045 14643 27079
rect 14609 26977 14643 27011
rect 14609 26909 14643 26943
rect 14609 26841 14643 26875
rect 14609 26773 14643 26807
rect 14609 26705 14643 26739
rect 14609 26637 14643 26671
rect 14609 26569 14643 26603
rect 14609 26501 14643 26535
rect 14609 26433 14643 26467
rect 14609 26365 14643 26399
rect 14609 26297 14643 26331
rect 14609 26229 14643 26263
rect 14609 26161 14643 26195
rect 14609 26093 14643 26127
rect 14609 26025 14643 26059
rect 14609 25957 14643 25991
rect 14609 25889 14643 25923
rect 14609 25821 14643 25855
rect 14609 25753 14643 25787
rect 14609 25685 14643 25719
rect 14609 25617 14643 25651
rect 14609 25549 14643 25583
rect 14609 25481 14643 25515
rect 14609 25413 14643 25447
rect 14609 25345 14643 25379
rect 14609 25277 14643 25311
rect 14609 25209 14643 25243
rect 14609 25141 14643 25175
rect 14609 25073 14643 25107
rect 14609 25005 14643 25039
rect 14609 24937 14643 24971
rect 14609 24869 14643 24903
rect 14609 24801 14643 24835
rect 14609 24733 14643 24767
rect 14609 24665 14643 24699
rect 14609 24597 14643 24631
rect 14609 24529 14643 24563
rect 14609 24461 14643 24495
rect 14609 24393 14643 24427
rect 14609 24325 14643 24359
rect 14609 24257 14643 24291
rect 14609 24189 14643 24223
rect 14609 24121 14643 24155
rect 14609 24053 14643 24087
rect 14609 23985 14643 24019
rect 14609 23917 14643 23951
rect 14609 23849 14643 23883
rect 14609 23781 14643 23815
rect 14609 23713 14643 23747
rect 14609 23645 14643 23679
rect 14609 23577 14643 23611
rect 14609 23509 14643 23543
rect 14609 23441 14643 23475
rect 14609 23373 14643 23407
rect 14609 23305 14643 23339
rect 14609 23237 14643 23271
rect 14609 23169 14643 23203
rect 14609 23101 14643 23135
rect 14609 23033 14643 23067
rect 14609 22965 14643 22999
rect 14609 22897 14643 22931
rect 14609 22829 14643 22863
rect 14609 22761 14643 22795
rect 14609 22693 14643 22727
rect 14609 22625 14643 22659
rect 14609 22557 14643 22591
rect 14609 22489 14643 22523
rect 14609 22421 14643 22455
rect 14609 22353 14643 22387
rect 14609 22285 14643 22319
rect 14609 22217 14643 22251
rect 14609 22149 14643 22183
rect 14609 22081 14643 22115
rect 14609 22013 14643 22047
rect 14609 21945 14643 21979
rect 14609 21877 14643 21911
rect 14609 21809 14643 21843
rect 14609 21741 14643 21775
rect 14609 21673 14643 21707
rect 14609 21605 14643 21639
rect 14609 21537 14643 21571
rect 14609 21469 14643 21503
rect 14609 21401 14643 21435
rect 14609 21333 14643 21367
rect 14609 21265 14643 21299
rect 14609 21197 14643 21231
rect 14609 21129 14643 21163
rect 14609 21061 14643 21095
rect 14609 20993 14643 21027
rect 14609 20925 14643 20959
rect 14609 20857 14643 20891
rect 14609 20789 14643 20823
rect 14609 20721 14643 20755
rect 14609 20653 14643 20687
rect 14609 20585 14643 20619
rect 14609 20517 14643 20551
rect 14609 20449 14643 20483
rect 14609 20381 14643 20415
rect 14609 20313 14643 20347
rect 14609 20245 14643 20279
rect 14609 20177 14643 20211
rect 14609 20109 14643 20143
rect 14609 20041 14643 20075
rect 14609 19973 14643 20007
rect 14609 19905 14643 19939
rect 14609 19837 14643 19871
rect 14609 19769 14643 19803
rect 14609 19701 14643 19735
rect 14609 19633 14643 19667
rect 14609 19565 14643 19599
rect 14609 19497 14643 19531
rect 14609 19429 14643 19463
rect 14609 19361 14643 19395
rect 14609 19293 14643 19327
rect 14609 19225 14643 19259
rect 14609 19157 14643 19191
rect 14609 19089 14643 19123
rect 14609 19021 14643 19055
rect 14609 18953 14643 18987
rect 14609 18885 14643 18919
rect 14609 18817 14643 18851
rect 14609 18749 14643 18783
rect 14609 18681 14643 18715
rect 14609 18613 14643 18647
rect 14609 18545 14643 18579
rect 14609 18477 14643 18511
rect 14609 18409 14643 18443
rect 14609 18341 14643 18375
rect 14609 18273 14643 18307
rect 14609 18205 14643 18239
rect 14609 18137 14643 18171
rect 14609 18069 14643 18103
rect 14609 18001 14643 18035
rect 14609 17933 14643 17967
rect 14609 17865 14643 17899
rect 14609 17797 14643 17831
rect 14609 17729 14643 17763
rect 14609 17661 14643 17695
rect 14609 17593 14643 17627
rect 14609 17525 14643 17559
rect 14609 17457 14643 17491
rect 14609 17389 14643 17423
rect 14609 17321 14643 17355
rect 14609 17253 14643 17287
rect 14609 17185 14643 17219
rect 14609 17117 14643 17151
rect 14609 17049 14643 17083
rect 14609 16981 14643 17015
rect 14609 16913 14643 16947
rect 14609 16845 14643 16879
rect 14609 16777 14643 16811
rect 14609 16709 14643 16743
rect 14609 16641 14643 16675
rect 14609 16573 14643 16607
rect 14609 16505 14643 16539
rect 14609 16437 14643 16471
rect 14609 16369 14643 16403
rect 14609 16301 14643 16335
rect 14609 16233 14643 16267
rect 14609 16165 14643 16199
rect 14609 16097 14643 16131
rect 14609 16029 14643 16063
rect 14609 15961 14643 15995
rect 14609 15893 14643 15927
rect 14609 15825 14643 15859
rect 14609 15757 14643 15791
rect 14609 15689 14643 15723
rect 14609 15621 14643 15655
rect 14609 15553 14643 15587
rect 14609 15485 14643 15519
rect 14609 15417 14643 15451
rect 14609 15349 14643 15383
rect 14609 15281 14643 15315
rect 14609 15213 14643 15247
rect 14609 15145 14643 15179
rect 14609 15077 14643 15111
rect 14609 15009 14643 15043
rect 14609 14941 14643 14975
rect 14609 14873 14643 14907
rect 14609 14805 14643 14839
rect 14609 14737 14643 14771
rect 14609 14669 14643 14703
rect 14609 14601 14643 14635
rect 14609 14533 14643 14567
rect 14609 14465 14643 14499
rect 14609 14397 14643 14431
rect 14609 14329 14643 14363
rect 14609 14261 14643 14295
rect 14609 14193 14643 14227
rect 14609 14125 14643 14159
rect 14609 14057 14643 14091
rect 14609 13989 14643 14023
rect 14609 13921 14643 13955
rect 14609 13853 14643 13887
rect 14609 13785 14643 13819
rect 14609 13717 14643 13751
rect 14609 13649 14643 13683
rect 14609 13581 14643 13615
rect 14609 13513 14643 13547
rect 14609 13445 14643 13479
rect 14609 13377 14643 13411
rect 14609 13309 14643 13343
rect 14609 13241 14643 13275
rect 14609 13173 14643 13207
rect 14609 13105 14643 13139
rect 14609 13037 14643 13071
rect 14609 12969 14643 13003
rect 14609 12901 14643 12935
rect 14609 12833 14643 12867
rect 14609 12765 14643 12799
rect 14609 12697 14643 12731
rect 14609 12629 14643 12663
rect 14609 12561 14643 12595
rect 14609 12493 14643 12527
rect 14609 12425 14643 12459
rect 14609 12357 14643 12391
rect 14609 12289 14643 12323
rect 14609 12221 14643 12255
rect 14609 12153 14643 12187
rect 14609 12085 14643 12119
rect 14609 12017 14643 12051
rect 14609 11949 14643 11983
rect 14609 11881 14643 11915
rect 14609 11813 14643 11847
rect 14609 11745 14643 11779
rect 14609 11677 14643 11711
rect 14609 11609 14643 11643
rect 14609 11541 14643 11575
rect 14609 11473 14643 11507
rect 14609 11405 14643 11439
rect 14609 11337 14643 11371
rect 14609 11269 14643 11303
rect 14609 11201 14643 11235
rect 14609 11133 14643 11167
rect 14609 11065 14643 11099
rect 14609 10997 14643 11031
rect 14609 10929 14643 10963
rect 14609 10861 14643 10895
rect 14609 10793 14643 10827
rect 14609 10725 14643 10759
rect 14609 10657 14643 10691
rect 14609 10589 14643 10623
rect 14609 10521 14643 10555
rect 14609 10453 14643 10487
rect 14609 10385 14643 10419
rect 14609 10317 14643 10351
rect 14609 10249 14643 10283
rect 14609 10181 14643 10215
rect 14609 10113 14643 10147
rect 14609 10045 14643 10079
rect 14609 9977 14643 10011
rect 14609 9909 14643 9943
rect 14609 9841 14643 9875
rect 14609 9773 14643 9807
rect 14609 9705 14643 9739
rect 322 9645 356 9679
rect 322 9577 356 9611
rect 14609 9637 14643 9671
rect 14609 9569 14643 9603
rect 510 9420 544 9454
rect 578 9420 612 9454
rect 646 9420 680 9454
rect 714 9420 748 9454
rect 782 9420 816 9454
rect 850 9420 884 9454
rect 918 9420 952 9454
rect 986 9420 1020 9454
rect 1054 9420 1088 9454
rect 1122 9420 1156 9454
rect 1190 9420 1224 9454
rect 1258 9420 1292 9454
rect 1326 9420 1360 9454
rect 1394 9420 1428 9454
rect 1462 9420 1496 9454
rect 1530 9420 1564 9454
rect 1598 9420 1632 9454
rect 1666 9420 1700 9454
rect 1734 9420 1768 9454
rect 1802 9420 1836 9454
rect 1870 9420 1904 9454
rect 1938 9420 1972 9454
rect 2006 9420 2040 9454
rect 2074 9420 2108 9454
rect 2142 9420 2176 9454
rect 2210 9420 2244 9454
rect 2278 9420 2312 9454
rect 2346 9420 2380 9454
rect 2414 9420 2448 9454
rect 2482 9420 2516 9454
rect 2550 9420 2584 9454
rect 2618 9420 2652 9454
rect 2686 9420 2720 9454
rect 2754 9420 2788 9454
rect 2822 9420 2856 9454
rect 2890 9420 2924 9454
rect 2958 9420 2992 9454
rect 3026 9420 3060 9454
rect 3094 9420 3128 9454
rect 3162 9420 3196 9454
rect 3230 9420 3264 9454
rect 3298 9420 3332 9454
rect 3366 9420 3400 9454
rect 3434 9420 3468 9454
rect 3502 9420 3536 9454
rect 3570 9420 3604 9454
rect 3638 9420 3672 9454
rect 3706 9420 3740 9454
rect 3774 9420 3808 9454
rect 3842 9420 3876 9454
rect 3910 9420 3944 9454
rect 3978 9420 4012 9454
rect 4046 9420 4080 9454
rect 4114 9420 4148 9454
rect 4182 9420 4216 9454
rect 4250 9420 4284 9454
rect 4318 9420 4352 9454
rect 4386 9420 4420 9454
rect 4454 9420 4488 9454
rect 4522 9420 4556 9454
rect 4590 9420 4624 9454
rect 4658 9420 4692 9454
rect 4726 9420 4760 9454
rect 4794 9420 4828 9454
rect 4862 9420 4896 9454
rect 4930 9420 4964 9454
rect 4998 9420 5032 9454
rect 5066 9420 5100 9454
rect 5134 9420 5168 9454
rect 5202 9420 5236 9454
rect 5270 9420 5304 9454
rect 5338 9420 5372 9454
rect 5406 9420 5440 9454
rect 5474 9420 5508 9454
rect 5542 9420 5576 9454
rect 5610 9420 5644 9454
rect 5678 9420 5712 9454
rect 5746 9420 5780 9454
rect 5814 9420 5848 9454
rect 5882 9420 5916 9454
rect 5950 9420 5984 9454
rect 6018 9420 6052 9454
rect 6086 9420 6120 9454
rect 6154 9420 6188 9454
rect 6222 9420 6256 9454
rect 6290 9420 6324 9454
rect 6358 9420 6392 9454
rect 6426 9420 6460 9454
rect 6494 9420 6528 9454
rect 6562 9420 6596 9454
rect 6630 9420 6664 9454
rect 6698 9420 6732 9454
rect 6766 9420 6800 9454
rect 6834 9420 6868 9454
rect 6902 9420 6936 9454
rect 6970 9420 7004 9454
rect 7038 9420 7072 9454
rect 7106 9420 7140 9454
rect 7174 9420 7208 9454
rect 7242 9420 7276 9454
rect 7310 9420 7344 9454
rect 7378 9420 7412 9454
rect 7446 9420 7480 9454
rect 7514 9420 7548 9454
rect 7582 9420 7616 9454
rect 7650 9420 7684 9454
rect 7718 9420 7752 9454
rect 7786 9420 7820 9454
rect 7854 9420 7888 9454
rect 7922 9420 7956 9454
rect 7990 9420 8024 9454
rect 8058 9420 8092 9454
rect 8126 9420 8160 9454
rect 8194 9420 8228 9454
rect 8262 9420 8296 9454
rect 8330 9420 8364 9454
rect 8398 9420 8432 9454
rect 8466 9420 8500 9454
rect 8534 9420 8568 9454
rect 8602 9420 8636 9454
rect 8670 9420 8704 9454
rect 8738 9420 8772 9454
rect 8806 9420 8840 9454
rect 8874 9420 8908 9454
rect 8942 9420 8976 9454
rect 9010 9420 9044 9454
rect 9078 9420 9112 9454
rect 9146 9420 9180 9454
rect 9214 9420 9248 9454
rect 9282 9420 9316 9454
rect 9350 9420 9384 9454
rect 9418 9420 9452 9454
rect 9486 9420 9520 9454
rect 9554 9420 9588 9454
rect 9622 9420 9656 9454
rect 9690 9420 9724 9454
rect 9758 9420 9792 9454
rect 9826 9420 9860 9454
rect 9894 9420 9928 9454
rect 9962 9420 9996 9454
rect 10030 9420 10064 9454
rect 10098 9420 10132 9454
rect 10166 9420 10200 9454
rect 10234 9420 10268 9454
rect 10302 9420 10336 9454
rect 10370 9420 10404 9454
rect 10438 9420 10472 9454
rect 10506 9420 10540 9454
rect 10574 9420 10608 9454
rect 10642 9420 10676 9454
rect 10710 9420 10744 9454
rect 10778 9420 10812 9454
rect 10846 9420 10880 9454
rect 10914 9420 10948 9454
rect 10982 9420 11016 9454
rect 11050 9420 11084 9454
rect 11118 9420 11152 9454
rect 11186 9420 11220 9454
rect 11254 9420 11288 9454
rect 11322 9420 11356 9454
rect 11390 9420 11424 9454
rect 11458 9420 11492 9454
rect 11526 9420 11560 9454
rect 11594 9420 11628 9454
rect 11662 9420 11696 9454
rect 11730 9420 11764 9454
rect 11798 9420 11832 9454
rect 11866 9420 11900 9454
rect 11934 9420 11968 9454
rect 12002 9420 12036 9454
rect 12070 9420 12104 9454
rect 12138 9420 12172 9454
rect 12206 9420 12240 9454
rect 12274 9420 12308 9454
rect 12342 9420 12376 9454
rect 12410 9420 12444 9454
rect 12478 9420 12512 9454
rect 12546 9420 12580 9454
rect 12614 9420 12648 9454
rect 12682 9420 12716 9454
rect 12750 9420 12784 9454
rect 12818 9420 12852 9454
rect 12886 9420 12920 9454
rect 12954 9420 12988 9454
rect 13022 9420 13056 9454
rect 13090 9420 13124 9454
rect 13158 9420 13192 9454
rect 13226 9420 13260 9454
rect 13294 9420 13328 9454
rect 13362 9420 13396 9454
rect 13430 9420 13464 9454
rect 13498 9420 13532 9454
rect 13566 9420 13600 9454
rect 13634 9420 13668 9454
rect 13702 9420 13736 9454
rect 13770 9420 13804 9454
rect 13838 9420 13872 9454
rect 13906 9420 13940 9454
rect 13974 9420 14008 9454
rect 14042 9420 14076 9454
rect 14110 9420 14144 9454
rect 14178 9420 14212 9454
rect 14246 9420 14280 9454
rect 14314 9420 14348 9454
rect 14382 9420 14416 9454
rect 14450 9420 14484 9454
<< mvnsubdiffcont >>
rect 773 36143 807 36177
rect 841 36143 875 36177
rect 909 36143 943 36177
rect 977 36143 1011 36177
rect 1045 36143 1079 36177
rect 1113 36143 1147 36177
rect 1181 36143 1215 36177
rect 1249 36143 1283 36177
rect 1317 36143 1351 36177
rect 1385 36143 1419 36177
rect 1453 36143 1487 36177
rect 1521 36143 1555 36177
rect 1589 36143 1623 36177
rect 1657 36143 1691 36177
rect 1725 36143 1759 36177
rect 1793 36143 1827 36177
rect 1861 36143 1895 36177
rect 1929 36143 1963 36177
rect 1997 36143 2031 36177
rect 2065 36143 2099 36177
rect 2133 36143 2167 36177
rect 2201 36143 2235 36177
rect 2269 36143 2303 36177
rect 2337 36143 2371 36177
rect 2405 36143 2439 36177
rect 2473 36143 2507 36177
rect 2541 36143 2575 36177
rect 2609 36143 2643 36177
rect 2677 36143 2711 36177
rect 2745 36143 2779 36177
rect 2813 36143 2847 36177
rect 2881 36143 2915 36177
rect 2949 36143 2983 36177
rect 3017 36143 3051 36177
rect 3085 36143 3119 36177
rect 3153 36143 3187 36177
rect 3221 36143 3255 36177
rect 3289 36143 3323 36177
rect 3357 36143 3391 36177
rect 3425 36143 3459 36177
rect 3493 36143 3527 36177
rect 3561 36143 3595 36177
rect 3629 36143 3663 36177
rect 3697 36143 3731 36177
rect 3765 36143 3799 36177
rect 3833 36143 3867 36177
rect 3901 36143 3935 36177
rect 3969 36143 4003 36177
rect 4037 36143 4071 36177
rect 4105 36143 4139 36177
rect 4173 36143 4207 36177
rect 4241 36143 4275 36177
rect 4309 36143 4343 36177
rect 4377 36143 4411 36177
rect 4445 36143 4479 36177
rect 4513 36143 4547 36177
rect 4581 36143 4615 36177
rect 4649 36143 4683 36177
rect 4717 36143 4751 36177
rect 4785 36143 4819 36177
rect 4853 36143 4887 36177
rect 4921 36143 4955 36177
rect 4989 36143 5023 36177
rect 5057 36143 5091 36177
rect 5125 36143 5159 36177
rect 5193 36143 5227 36177
rect 5261 36143 5295 36177
rect 5329 36143 5363 36177
rect 5397 36143 5431 36177
rect 5465 36143 5499 36177
rect 5533 36143 5567 36177
rect 5601 36143 5635 36177
rect 5669 36143 5703 36177
rect 5737 36143 5771 36177
rect 5805 36143 5839 36177
rect 5873 36143 5907 36177
rect 5941 36143 5975 36177
rect 6009 36143 6043 36177
rect 6077 36143 6111 36177
rect 6145 36143 6179 36177
rect 6213 36143 6247 36177
rect 6281 36143 6315 36177
rect 6349 36143 6383 36177
rect 6417 36143 6451 36177
rect 6485 36143 6519 36177
rect 6553 36143 6587 36177
rect 6621 36143 6655 36177
rect 6689 36143 6723 36177
rect 6757 36143 6791 36177
rect 6825 36143 6859 36177
rect 6893 36143 6927 36177
rect 6961 36143 6995 36177
rect 7029 36143 7063 36177
rect 7097 36143 7131 36177
rect 7165 36143 7199 36177
rect 7233 36143 7267 36177
rect 7301 36143 7335 36177
rect 7369 36143 7403 36177
rect 7437 36143 7471 36177
rect 7505 36143 7539 36177
rect 7573 36143 7607 36177
rect 7641 36143 7675 36177
rect 7709 36143 7743 36177
rect 7777 36143 7811 36177
rect 7845 36143 7879 36177
rect 7913 36143 7947 36177
rect 7981 36143 8015 36177
rect 8049 36143 8083 36177
rect 8117 36143 8151 36177
rect 8185 36143 8219 36177
rect 8253 36143 8287 36177
rect 8321 36143 8355 36177
rect 8389 36143 8423 36177
rect 8457 36143 8491 36177
rect 8525 36143 8559 36177
rect 8593 36143 8627 36177
rect 8661 36143 8695 36177
rect 8729 36143 8763 36177
rect 8797 36143 8831 36177
rect 8865 36143 8899 36177
rect 8933 36143 8967 36177
rect 9001 36143 9035 36177
rect 9069 36143 9103 36177
rect 9137 36143 9171 36177
rect 9205 36143 9239 36177
rect 9273 36143 9307 36177
rect 9341 36143 9375 36177
rect 9409 36143 9443 36177
rect 9477 36143 9511 36177
rect 9545 36143 9579 36177
rect 9613 36143 9647 36177
rect 9681 36143 9715 36177
rect 9749 36143 9783 36177
rect 9817 36143 9851 36177
rect 9885 36143 9919 36177
rect 9953 36143 9987 36177
rect 10021 36143 10055 36177
rect 10089 36143 10123 36177
rect 10157 36143 10191 36177
rect 10225 36143 10259 36177
rect 10293 36143 10327 36177
rect 10361 36143 10395 36177
rect 10429 36143 10463 36177
rect 10497 36143 10531 36177
rect 10565 36143 10599 36177
rect 10633 36143 10667 36177
rect 10701 36143 10735 36177
rect 10769 36143 10803 36177
rect 10837 36143 10871 36177
rect 10905 36143 10939 36177
rect 10973 36143 11007 36177
rect 11041 36143 11075 36177
rect 11109 36143 11143 36177
rect 11177 36143 11211 36177
rect 11245 36143 11279 36177
rect 11313 36143 11347 36177
rect 11381 36143 11415 36177
rect 11449 36143 11483 36177
rect 11517 36143 11551 36177
rect 11585 36143 11619 36177
rect 11653 36143 11687 36177
rect 11721 36143 11755 36177
rect 11789 36143 11823 36177
rect 11857 36143 11891 36177
rect 11925 36143 11959 36177
rect 11993 36143 12027 36177
rect 12061 36143 12095 36177
rect 12129 36143 12163 36177
rect 12197 36143 12231 36177
rect 12265 36143 12299 36177
rect 12333 36143 12367 36177
rect 12401 36143 12435 36177
rect 12469 36143 12503 36177
rect 12537 36143 12571 36177
rect 12605 36143 12639 36177
rect 12673 36143 12707 36177
rect 12741 36143 12775 36177
rect 12809 36143 12843 36177
rect 12877 36143 12911 36177
rect 12945 36143 12979 36177
rect 13013 36143 13047 36177
rect 13081 36143 13115 36177
rect 13149 36143 13183 36177
rect 13217 36143 13251 36177
rect 13285 36143 13319 36177
rect 13353 36143 13387 36177
rect 13421 36143 13455 36177
rect 13489 36143 13523 36177
rect 13557 36143 13591 36177
rect 13625 36143 13659 36177
rect 13693 36143 13727 36177
rect 13761 36143 13795 36177
rect 13829 36143 13863 36177
rect 13897 36143 13931 36177
rect 13965 36143 13999 36177
rect 14033 36143 14067 36177
rect 14101 36143 14135 36177
rect 14169 36143 14203 36177
rect 646 35998 680 36032
rect 646 35930 680 35964
rect 646 35862 680 35896
rect 646 35794 680 35828
rect 646 35726 680 35760
rect 646 35658 680 35692
rect 646 35590 680 35624
rect 646 35522 680 35556
rect 646 35454 680 35488
rect 646 35386 680 35420
rect 646 35318 680 35352
rect 646 35250 680 35284
rect 646 35182 680 35216
rect 646 35114 680 35148
rect 646 35046 680 35080
rect 646 34978 680 35012
rect 646 34910 680 34944
rect 646 34842 680 34876
rect 646 34774 680 34808
rect 646 34706 680 34740
rect 14297 35998 14331 36032
rect 14297 35930 14331 35964
rect 14297 35862 14331 35896
rect 14297 35794 14331 35828
rect 14297 35726 14331 35760
rect 14297 35658 14331 35692
rect 14297 35590 14331 35624
rect 14297 35522 14331 35556
rect 14297 35454 14331 35488
rect 14297 35386 14331 35420
rect 14297 35318 14331 35352
rect 14297 35250 14331 35284
rect 14297 35182 14331 35216
rect 14297 35114 14331 35148
rect 14297 35046 14331 35080
rect 14297 34978 14331 35012
rect 14297 34910 14331 34944
rect 14297 34842 14331 34876
rect 14297 34774 14331 34808
rect 14297 34706 14331 34740
rect 646 34638 680 34672
rect 646 34570 680 34604
rect 646 34502 680 34536
rect 646 34434 680 34468
rect 646 34366 680 34400
rect 646 34298 680 34332
rect 646 34230 680 34264
rect 646 34162 680 34196
rect 646 34094 680 34128
rect 646 34026 680 34060
rect 646 33958 680 33992
rect 646 33890 680 33924
rect 646 33822 680 33856
rect 646 33754 680 33788
rect 646 33686 680 33720
rect 646 33618 680 33652
rect 646 33550 680 33584
rect 646 33482 680 33516
rect 646 33414 680 33448
rect 646 33346 680 33380
rect 646 33278 680 33312
rect 646 33210 680 33244
rect 646 33142 680 33176
rect 646 33074 680 33108
rect 646 33006 680 33040
rect 646 32938 680 32972
rect 646 32870 680 32904
rect 646 32802 680 32836
rect 646 32734 680 32768
rect 646 32666 680 32700
rect 646 32598 680 32632
rect 646 32530 680 32564
rect 646 32462 680 32496
rect 646 32394 680 32428
rect 646 32326 680 32360
rect 646 32258 680 32292
rect 646 32190 680 32224
rect 646 32122 680 32156
rect 646 32054 680 32088
rect 646 31986 680 32020
rect 646 31918 680 31952
rect 646 31850 680 31884
rect 646 31782 680 31816
rect 646 31714 680 31748
rect 646 31646 680 31680
rect 646 31578 680 31612
rect 646 31510 680 31544
rect 646 31442 680 31476
rect 646 31374 680 31408
rect 646 31306 680 31340
rect 646 31238 680 31272
rect 646 31170 680 31204
rect 646 31102 680 31136
rect 646 31034 680 31068
rect 646 30966 680 31000
rect 646 30898 680 30932
rect 646 30830 680 30864
rect 646 30762 680 30796
rect 646 30694 680 30728
rect 646 30626 680 30660
rect 646 30558 680 30592
rect 646 30490 680 30524
rect 646 30422 680 30456
rect 646 30354 680 30388
rect 646 30286 680 30320
rect 646 30218 680 30252
rect 646 30150 680 30184
rect 646 30082 680 30116
rect 646 30014 680 30048
rect 646 29946 680 29980
rect 646 29878 680 29912
rect 646 29810 680 29844
rect 646 29742 680 29776
rect 646 29674 680 29708
rect 646 29606 680 29640
rect 646 29538 680 29572
rect 646 29470 680 29504
rect 646 29402 680 29436
rect 646 29334 680 29368
rect 646 29266 680 29300
rect 646 29198 680 29232
rect 646 29130 680 29164
rect 646 29062 680 29096
rect 646 28994 680 29028
rect 646 28926 680 28960
rect 646 28858 680 28892
rect 646 28790 680 28824
rect 646 28722 680 28756
rect 646 28654 680 28688
rect 646 28586 680 28620
rect 646 28518 680 28552
rect 646 28450 680 28484
rect 646 28382 680 28416
rect 646 28314 680 28348
rect 646 28246 680 28280
rect 646 28178 680 28212
rect 646 28110 680 28144
rect 646 28042 680 28076
rect 646 27974 680 28008
rect 646 27906 680 27940
rect 646 27838 680 27872
rect 646 27770 680 27804
rect 646 27702 680 27736
rect 646 27634 680 27668
rect 646 27566 680 27600
rect 646 27498 680 27532
rect 646 27430 680 27464
rect 646 27362 680 27396
rect 646 27294 680 27328
rect 646 27226 680 27260
rect 646 27158 680 27192
rect 646 27090 680 27124
rect 646 27022 680 27056
rect 646 26954 680 26988
rect 646 26886 680 26920
rect 646 26818 680 26852
rect 646 26750 680 26784
rect 646 26682 680 26716
rect 646 26614 680 26648
rect 646 26546 680 26580
rect 646 26478 680 26512
rect 646 26410 680 26444
rect 646 26342 680 26376
rect 646 26274 680 26308
rect 646 26206 680 26240
rect 646 26138 680 26172
rect 646 26070 680 26104
rect 646 26002 680 26036
rect 646 25934 680 25968
rect 646 25866 680 25900
rect 646 25798 680 25832
rect 646 25730 680 25764
rect 646 25662 680 25696
rect 646 25594 680 25628
rect 646 25526 680 25560
rect 646 25458 680 25492
rect 646 25390 680 25424
rect 646 25322 680 25356
rect 646 25254 680 25288
rect 646 25186 680 25220
rect 646 25118 680 25152
rect 646 25050 680 25084
rect 646 24982 680 25016
rect 646 24914 680 24948
rect 646 24846 680 24880
rect 646 24778 680 24812
rect 646 24710 680 24744
rect 646 24642 680 24676
rect 646 24574 680 24608
rect 646 24506 680 24540
rect 646 24438 680 24472
rect 646 24370 680 24404
rect 646 24302 680 24336
rect 646 24234 680 24268
rect 646 24166 680 24200
rect 646 24098 680 24132
rect 646 24030 680 24064
rect 646 23962 680 23996
rect 646 23894 680 23928
rect 646 23826 680 23860
rect 646 23758 680 23792
rect 646 23690 680 23724
rect 646 23622 680 23656
rect 646 23554 680 23588
rect 646 23486 680 23520
rect 646 23418 680 23452
rect 646 23350 680 23384
rect 646 23282 680 23316
rect 646 23214 680 23248
rect 646 23146 680 23180
rect 646 23078 680 23112
rect 646 23010 680 23044
rect 646 22942 680 22976
rect 646 22874 680 22908
rect 646 22806 680 22840
rect 646 22738 680 22772
rect 646 22670 680 22704
rect 646 22602 680 22636
rect 646 22534 680 22568
rect 646 22466 680 22500
rect 646 22398 680 22432
rect 646 22330 680 22364
rect 646 22262 680 22296
rect 646 22194 680 22228
rect 646 22126 680 22160
rect 646 22058 680 22092
rect 646 21990 680 22024
rect 646 21922 680 21956
rect 646 21854 680 21888
rect 646 21786 680 21820
rect 646 21718 680 21752
rect 646 21650 680 21684
rect 646 21582 680 21616
rect 646 21514 680 21548
rect 646 21446 680 21480
rect 646 21378 680 21412
rect 646 21310 680 21344
rect 646 21242 680 21276
rect 646 21174 680 21208
rect 646 21106 680 21140
rect 646 21038 680 21072
rect 646 20970 680 21004
rect 646 20902 680 20936
rect 646 20834 680 20868
rect 646 20766 680 20800
rect 646 20698 680 20732
rect 646 20630 680 20664
rect 646 20562 680 20596
rect 646 20494 680 20528
rect 646 20426 680 20460
rect 646 20358 680 20392
rect 646 20290 680 20324
rect 646 20222 680 20256
rect 646 20154 680 20188
rect 646 20086 680 20120
rect 646 20018 680 20052
rect 646 19950 680 19984
rect 646 19882 680 19916
rect 646 19814 680 19848
rect 646 19746 680 19780
rect 646 19678 680 19712
rect 646 19610 680 19644
rect 646 19542 680 19576
rect 646 19474 680 19508
rect 646 19406 680 19440
rect 646 19338 680 19372
rect 646 19270 680 19304
rect 646 19202 680 19236
rect 646 19134 680 19168
rect 646 19066 680 19100
rect 646 18998 680 19032
rect 646 18930 680 18964
rect 646 18862 680 18896
rect 646 18794 680 18828
rect 646 18726 680 18760
rect 646 18658 680 18692
rect 646 18590 680 18624
rect 646 18522 680 18556
rect 646 18454 680 18488
rect 646 18386 680 18420
rect 646 18318 680 18352
rect 646 18250 680 18284
rect 646 18182 680 18216
rect 646 18114 680 18148
rect 646 18046 680 18080
rect 646 17978 680 18012
rect 646 17910 680 17944
rect 646 17842 680 17876
rect 646 17774 680 17808
rect 646 17706 680 17740
rect 646 17638 680 17672
rect 646 17570 680 17604
rect 646 17502 680 17536
rect 646 17434 680 17468
rect 646 17366 680 17400
rect 646 17298 680 17332
rect 646 17230 680 17264
rect 646 17162 680 17196
rect 646 17094 680 17128
rect 646 17026 680 17060
rect 646 16958 680 16992
rect 646 16890 680 16924
rect 646 16822 680 16856
rect 646 16754 680 16788
rect 646 16686 680 16720
rect 646 16618 680 16652
rect 646 16550 680 16584
rect 646 16482 680 16516
rect 646 16414 680 16448
rect 646 16346 680 16380
rect 646 16278 680 16312
rect 646 16210 680 16244
rect 646 16142 680 16176
rect 646 16074 680 16108
rect 646 16006 680 16040
rect 646 15938 680 15972
rect 646 15870 680 15904
rect 646 15802 680 15836
rect 646 15734 680 15768
rect 646 15666 680 15700
rect 646 15598 680 15632
rect 646 15530 680 15564
rect 646 15462 680 15496
rect 646 15394 680 15428
rect 646 15326 680 15360
rect 646 15258 680 15292
rect 646 15190 680 15224
rect 646 15122 680 15156
rect 646 15054 680 15088
rect 646 14986 680 15020
rect 646 14918 680 14952
rect 646 14850 680 14884
rect 646 14782 680 14816
rect 646 14714 680 14748
rect 646 14646 680 14680
rect 646 14578 680 14612
rect 646 14510 680 14544
rect 646 14442 680 14476
rect 646 14374 680 14408
rect 646 14306 680 14340
rect 646 14238 680 14272
rect 646 14170 680 14204
rect 646 14102 680 14136
rect 646 14034 680 14068
rect 646 13966 680 14000
rect 646 13898 680 13932
rect 646 13830 680 13864
rect 646 13762 680 13796
rect 646 13694 680 13728
rect 646 13626 680 13660
rect 646 13558 680 13592
rect 646 13490 680 13524
rect 646 13422 680 13456
rect 646 13354 680 13388
rect 646 13286 680 13320
rect 646 13218 680 13252
rect 646 13150 680 13184
rect 646 13082 680 13116
rect 646 13014 680 13048
rect 646 12946 680 12980
rect 646 12878 680 12912
rect 646 12810 680 12844
rect 646 12742 680 12776
rect 646 12674 680 12708
rect 646 12606 680 12640
rect 646 12538 680 12572
rect 646 12470 680 12504
rect 646 12402 680 12436
rect 646 12334 680 12368
rect 646 12266 680 12300
rect 646 12198 680 12232
rect 646 12130 680 12164
rect 646 12062 680 12096
rect 646 11994 680 12028
rect 646 11926 680 11960
rect 646 11858 680 11892
rect 646 11790 680 11824
rect 646 11722 680 11756
rect 646 11654 680 11688
rect 646 11586 680 11620
rect 646 11518 680 11552
rect 646 11450 680 11484
rect 646 11382 680 11416
rect 646 11314 680 11348
rect 646 11246 680 11280
rect 646 11178 680 11212
rect 646 11110 680 11144
rect 646 11042 680 11076
rect 646 10974 680 11008
rect 646 10906 680 10940
rect 646 10838 680 10872
rect 646 10770 680 10804
rect 646 10702 680 10736
rect 646 10634 680 10668
rect 646 10566 680 10600
rect 646 10498 680 10532
rect 646 10430 680 10464
rect 646 10362 680 10396
rect 646 10294 680 10328
rect 646 10226 680 10260
rect 14297 34638 14331 34672
rect 14297 34570 14331 34604
rect 14297 34502 14331 34536
rect 14297 34434 14331 34468
rect 14297 34366 14331 34400
rect 14297 34298 14331 34332
rect 14297 34230 14331 34264
rect 14297 34162 14331 34196
rect 14297 34094 14331 34128
rect 14297 34026 14331 34060
rect 14297 33958 14331 33992
rect 14297 33890 14331 33924
rect 14297 33822 14331 33856
rect 14297 33754 14331 33788
rect 14297 33686 14331 33720
rect 14297 33618 14331 33652
rect 14297 33550 14331 33584
rect 14297 33482 14331 33516
rect 14297 33414 14331 33448
rect 14297 33346 14331 33380
rect 14297 33278 14331 33312
rect 14297 33210 14331 33244
rect 14297 33142 14331 33176
rect 14297 33074 14331 33108
rect 14297 33006 14331 33040
rect 14297 32938 14331 32972
rect 14297 32870 14331 32904
rect 14297 32802 14331 32836
rect 14297 32734 14331 32768
rect 14297 32666 14331 32700
rect 14297 32598 14331 32632
rect 14297 32530 14331 32564
rect 14297 32462 14331 32496
rect 14297 32394 14331 32428
rect 14297 32326 14331 32360
rect 14297 32258 14331 32292
rect 14297 32190 14331 32224
rect 14297 32122 14331 32156
rect 14297 32054 14331 32088
rect 14297 31986 14331 32020
rect 14297 31918 14331 31952
rect 14297 31850 14331 31884
rect 14297 31782 14331 31816
rect 14297 31714 14331 31748
rect 14297 31646 14331 31680
rect 14297 31578 14331 31612
rect 14297 31510 14331 31544
rect 14297 31442 14331 31476
rect 14297 31374 14331 31408
rect 14297 31306 14331 31340
rect 14297 31238 14331 31272
rect 14297 31170 14331 31204
rect 14297 31102 14331 31136
rect 14297 31034 14331 31068
rect 14297 30966 14331 31000
rect 14297 30898 14331 30932
rect 14297 30830 14331 30864
rect 14297 30762 14331 30796
rect 14297 30694 14331 30728
rect 14297 30626 14331 30660
rect 14297 30558 14331 30592
rect 14297 30490 14331 30524
rect 14297 30422 14331 30456
rect 14297 30354 14331 30388
rect 14297 30286 14331 30320
rect 14297 30218 14331 30252
rect 14297 30150 14331 30184
rect 14297 30082 14331 30116
rect 14297 30014 14331 30048
rect 14297 29946 14331 29980
rect 14297 29878 14331 29912
rect 14297 29810 14331 29844
rect 14297 29742 14331 29776
rect 14297 29674 14331 29708
rect 14297 29606 14331 29640
rect 14297 29538 14331 29572
rect 14297 29470 14331 29504
rect 14297 29402 14331 29436
rect 14297 29334 14331 29368
rect 14297 29266 14331 29300
rect 14297 29198 14331 29232
rect 14297 29130 14331 29164
rect 14297 29062 14331 29096
rect 14297 28994 14331 29028
rect 14297 28926 14331 28960
rect 14297 28858 14331 28892
rect 14297 28790 14331 28824
rect 14297 28722 14331 28756
rect 14297 28654 14331 28688
rect 14297 28586 14331 28620
rect 14297 28518 14331 28552
rect 14297 28450 14331 28484
rect 14297 28382 14331 28416
rect 14297 28314 14331 28348
rect 14297 28246 14331 28280
rect 14297 28178 14331 28212
rect 14297 28110 14331 28144
rect 14297 28042 14331 28076
rect 14297 27974 14331 28008
rect 14297 27906 14331 27940
rect 14297 27838 14331 27872
rect 14297 27770 14331 27804
rect 14297 27702 14331 27736
rect 14297 27634 14331 27668
rect 14297 27566 14331 27600
rect 14297 27498 14331 27532
rect 14297 27430 14331 27464
rect 14297 27362 14331 27396
rect 14297 27294 14331 27328
rect 14297 27226 14331 27260
rect 14297 27158 14331 27192
rect 14297 27090 14331 27124
rect 14297 27022 14331 27056
rect 14297 26954 14331 26988
rect 14297 26886 14331 26920
rect 14297 26818 14331 26852
rect 14297 26750 14331 26784
rect 14297 26682 14331 26716
rect 14297 26614 14331 26648
rect 14297 26546 14331 26580
rect 14297 26478 14331 26512
rect 14297 26410 14331 26444
rect 14297 26342 14331 26376
rect 14297 26274 14331 26308
rect 14297 26206 14331 26240
rect 14297 26138 14331 26172
rect 14297 26070 14331 26104
rect 14297 26002 14331 26036
rect 14297 25934 14331 25968
rect 14297 25866 14331 25900
rect 14297 25798 14331 25832
rect 14297 25730 14331 25764
rect 14297 25662 14331 25696
rect 14297 25594 14331 25628
rect 14297 25526 14331 25560
rect 14297 25458 14331 25492
rect 14297 25390 14331 25424
rect 14297 25322 14331 25356
rect 14297 25254 14331 25288
rect 14297 25186 14331 25220
rect 14297 25118 14331 25152
rect 14297 25050 14331 25084
rect 14297 24982 14331 25016
rect 14297 24914 14331 24948
rect 14297 24846 14331 24880
rect 14297 24778 14331 24812
rect 14297 24710 14331 24744
rect 14297 24642 14331 24676
rect 14297 24574 14331 24608
rect 14297 24506 14331 24540
rect 14297 24438 14331 24472
rect 14297 24370 14331 24404
rect 14297 24302 14331 24336
rect 14297 24234 14331 24268
rect 14297 24166 14331 24200
rect 14297 24098 14331 24132
rect 14297 24030 14331 24064
rect 14297 23962 14331 23996
rect 14297 23894 14331 23928
rect 14297 23826 14331 23860
rect 14297 23758 14331 23792
rect 14297 23690 14331 23724
rect 14297 23622 14331 23656
rect 14297 23554 14331 23588
rect 14297 23486 14331 23520
rect 14297 23418 14331 23452
rect 14297 23350 14331 23384
rect 14297 23282 14331 23316
rect 14297 23214 14331 23248
rect 14297 23146 14331 23180
rect 14297 23078 14331 23112
rect 14297 23010 14331 23044
rect 14297 22942 14331 22976
rect 14297 22874 14331 22908
rect 14297 22806 14331 22840
rect 14297 22738 14331 22772
rect 14297 22670 14331 22704
rect 14297 22602 14331 22636
rect 14297 22534 14331 22568
rect 14297 22466 14331 22500
rect 14297 22398 14331 22432
rect 14297 22330 14331 22364
rect 14297 22262 14331 22296
rect 14297 22194 14331 22228
rect 14297 22126 14331 22160
rect 14297 22058 14331 22092
rect 14297 21990 14331 22024
rect 14297 21922 14331 21956
rect 14297 21854 14331 21888
rect 14297 21786 14331 21820
rect 14297 21718 14331 21752
rect 14297 21650 14331 21684
rect 14297 21582 14331 21616
rect 14297 21514 14331 21548
rect 14297 21446 14331 21480
rect 14297 21378 14331 21412
rect 14297 21310 14331 21344
rect 14297 21242 14331 21276
rect 14297 21174 14331 21208
rect 14297 21106 14331 21140
rect 14297 21038 14331 21072
rect 14297 20970 14331 21004
rect 14297 20902 14331 20936
rect 14297 20834 14331 20868
rect 14297 20766 14331 20800
rect 14297 20698 14331 20732
rect 14297 20630 14331 20664
rect 14297 20562 14331 20596
rect 14297 20494 14331 20528
rect 14297 20426 14331 20460
rect 14297 20358 14331 20392
rect 14297 20290 14331 20324
rect 14297 20222 14331 20256
rect 14297 20154 14331 20188
rect 14297 20086 14331 20120
rect 14297 20018 14331 20052
rect 14297 19950 14331 19984
rect 14297 19882 14331 19916
rect 14297 19814 14331 19848
rect 14297 19746 14331 19780
rect 14297 19678 14331 19712
rect 14297 19610 14331 19644
rect 14297 19542 14331 19576
rect 14297 19474 14331 19508
rect 14297 19406 14331 19440
rect 14297 19338 14331 19372
rect 14297 19270 14331 19304
rect 14297 19202 14331 19236
rect 14297 19134 14331 19168
rect 14297 19066 14331 19100
rect 14297 18998 14331 19032
rect 14297 18930 14331 18964
rect 14297 18862 14331 18896
rect 14297 18794 14331 18828
rect 14297 18726 14331 18760
rect 14297 18658 14331 18692
rect 14297 18590 14331 18624
rect 14297 18522 14331 18556
rect 14297 18454 14331 18488
rect 14297 18386 14331 18420
rect 14297 18318 14331 18352
rect 14297 18250 14331 18284
rect 14297 18182 14331 18216
rect 14297 18114 14331 18148
rect 14297 18046 14331 18080
rect 14297 17978 14331 18012
rect 14297 17910 14331 17944
rect 14297 17842 14331 17876
rect 14297 17774 14331 17808
rect 14297 17706 14331 17740
rect 14297 17638 14331 17672
rect 14297 17570 14331 17604
rect 14297 17502 14331 17536
rect 14297 17434 14331 17468
rect 14297 17366 14331 17400
rect 14297 17298 14331 17332
rect 14297 17230 14331 17264
rect 14297 17162 14331 17196
rect 14297 17094 14331 17128
rect 14297 17026 14331 17060
rect 14297 16958 14331 16992
rect 14297 16890 14331 16924
rect 14297 16822 14331 16856
rect 14297 16754 14331 16788
rect 14297 16686 14331 16720
rect 14297 16618 14331 16652
rect 14297 16550 14331 16584
rect 14297 16482 14331 16516
rect 14297 16414 14331 16448
rect 14297 16346 14331 16380
rect 14297 16278 14331 16312
rect 14297 16210 14331 16244
rect 14297 16142 14331 16176
rect 14297 16074 14331 16108
rect 14297 16006 14331 16040
rect 14297 15938 14331 15972
rect 14297 15870 14331 15904
rect 14297 15802 14331 15836
rect 14297 15734 14331 15768
rect 14297 15666 14331 15700
rect 14297 15598 14331 15632
rect 14297 15530 14331 15564
rect 14297 15462 14331 15496
rect 14297 15394 14331 15428
rect 14297 15326 14331 15360
rect 14297 15258 14331 15292
rect 14297 15190 14331 15224
rect 14297 15122 14331 15156
rect 14297 15054 14331 15088
rect 14297 14986 14331 15020
rect 14297 14918 14331 14952
rect 14297 14850 14331 14884
rect 14297 14782 14331 14816
rect 14297 14714 14331 14748
rect 14297 14646 14331 14680
rect 14297 14578 14331 14612
rect 14297 14510 14331 14544
rect 14297 14442 14331 14476
rect 14297 14374 14331 14408
rect 14297 14306 14331 14340
rect 14297 14238 14331 14272
rect 14297 14170 14331 14204
rect 14297 14102 14331 14136
rect 14297 14034 14331 14068
rect 14297 13966 14331 14000
rect 14297 13898 14331 13932
rect 14297 13830 14331 13864
rect 14297 13762 14331 13796
rect 14297 13694 14331 13728
rect 14297 13626 14331 13660
rect 14297 13558 14331 13592
rect 14297 13490 14331 13524
rect 14297 13422 14331 13456
rect 14297 13354 14331 13388
rect 14297 13286 14331 13320
rect 14297 13218 14331 13252
rect 14297 13150 14331 13184
rect 14297 13082 14331 13116
rect 14297 13014 14331 13048
rect 14297 12946 14331 12980
rect 14297 12878 14331 12912
rect 14297 12810 14331 12844
rect 14297 12742 14331 12776
rect 14297 12674 14331 12708
rect 14297 12606 14331 12640
rect 14297 12538 14331 12572
rect 14297 12470 14331 12504
rect 14297 12402 14331 12436
rect 14297 12334 14331 12368
rect 14297 12266 14331 12300
rect 14297 12198 14331 12232
rect 14297 12130 14331 12164
rect 14297 12062 14331 12096
rect 14297 11994 14331 12028
rect 14297 11926 14331 11960
rect 14297 11858 14331 11892
rect 14297 11790 14331 11824
rect 14297 11722 14331 11756
rect 14297 11654 14331 11688
rect 14297 11586 14331 11620
rect 14297 11518 14331 11552
rect 14297 11450 14331 11484
rect 14297 11382 14331 11416
rect 14297 11314 14331 11348
rect 14297 11246 14331 11280
rect 14297 11178 14331 11212
rect 14297 11110 14331 11144
rect 14297 11042 14331 11076
rect 14297 10974 14331 11008
rect 14297 10906 14331 10940
rect 14297 10838 14331 10872
rect 14297 10770 14331 10804
rect 14297 10702 14331 10736
rect 14297 10634 14331 10668
rect 14297 10566 14331 10600
rect 14297 10498 14331 10532
rect 14297 10430 14331 10464
rect 14297 10362 14331 10396
rect 14297 10294 14331 10328
rect 14297 10226 14331 10260
rect 646 10158 680 10192
rect 646 10090 680 10124
rect 646 10022 680 10056
rect 646 9954 680 9988
rect 646 9886 680 9920
rect 14297 10158 14331 10192
rect 14297 10090 14331 10124
rect 14297 10022 14331 10056
rect 14297 9954 14331 9988
rect 14297 9886 14331 9920
rect 773 9741 807 9775
rect 841 9741 875 9775
rect 909 9741 943 9775
rect 977 9741 1011 9775
rect 1045 9741 1079 9775
rect 1113 9741 1147 9775
rect 1181 9741 1215 9775
rect 1249 9741 1283 9775
rect 1317 9741 1351 9775
rect 1385 9741 1419 9775
rect 1453 9741 1487 9775
rect 1521 9741 1555 9775
rect 1589 9741 1623 9775
rect 1657 9741 1691 9775
rect 1725 9741 1759 9775
rect 1793 9741 1827 9775
rect 1861 9741 1895 9775
rect 1929 9741 1963 9775
rect 1997 9741 2031 9775
rect 2065 9741 2099 9775
rect 2133 9741 2167 9775
rect 2201 9741 2235 9775
rect 2269 9741 2303 9775
rect 2337 9741 2371 9775
rect 2405 9741 2439 9775
rect 2473 9741 2507 9775
rect 2541 9741 2575 9775
rect 2609 9741 2643 9775
rect 2677 9741 2711 9775
rect 2745 9741 2779 9775
rect 2813 9741 2847 9775
rect 2881 9741 2915 9775
rect 2949 9741 2983 9775
rect 3017 9741 3051 9775
rect 3085 9741 3119 9775
rect 3153 9741 3187 9775
rect 3221 9741 3255 9775
rect 3289 9741 3323 9775
rect 3357 9741 3391 9775
rect 3425 9741 3459 9775
rect 3493 9741 3527 9775
rect 3561 9741 3595 9775
rect 3629 9741 3663 9775
rect 3697 9741 3731 9775
rect 3765 9741 3799 9775
rect 3833 9741 3867 9775
rect 3901 9741 3935 9775
rect 3969 9741 4003 9775
rect 4037 9741 4071 9775
rect 4105 9741 4139 9775
rect 4173 9741 4207 9775
rect 4241 9741 4275 9775
rect 4309 9741 4343 9775
rect 4377 9741 4411 9775
rect 4445 9741 4479 9775
rect 4513 9741 4547 9775
rect 4581 9741 4615 9775
rect 4649 9741 4683 9775
rect 4717 9741 4751 9775
rect 4785 9741 4819 9775
rect 4853 9741 4887 9775
rect 4921 9741 4955 9775
rect 4989 9741 5023 9775
rect 5057 9741 5091 9775
rect 5125 9741 5159 9775
rect 5193 9741 5227 9775
rect 5261 9741 5295 9775
rect 5329 9741 5363 9775
rect 5397 9741 5431 9775
rect 5465 9741 5499 9775
rect 5533 9741 5567 9775
rect 5601 9741 5635 9775
rect 5669 9741 5703 9775
rect 5737 9741 5771 9775
rect 5805 9741 5839 9775
rect 5873 9741 5907 9775
rect 5941 9741 5975 9775
rect 6009 9741 6043 9775
rect 6077 9741 6111 9775
rect 6145 9741 6179 9775
rect 6213 9741 6247 9775
rect 6281 9741 6315 9775
rect 6349 9741 6383 9775
rect 6417 9741 6451 9775
rect 6485 9741 6519 9775
rect 6553 9741 6587 9775
rect 6621 9741 6655 9775
rect 6689 9741 6723 9775
rect 6757 9741 6791 9775
rect 6825 9741 6859 9775
rect 6893 9741 6927 9775
rect 6961 9741 6995 9775
rect 7029 9741 7063 9775
rect 7097 9741 7131 9775
rect 7165 9741 7199 9775
rect 7233 9741 7267 9775
rect 7301 9741 7335 9775
rect 7369 9741 7403 9775
rect 7437 9741 7471 9775
rect 7505 9741 7539 9775
rect 7573 9741 7607 9775
rect 7641 9741 7675 9775
rect 7709 9741 7743 9775
rect 7777 9741 7811 9775
rect 7845 9741 7879 9775
rect 7913 9741 7947 9775
rect 7981 9741 8015 9775
rect 8049 9741 8083 9775
rect 8117 9741 8151 9775
rect 8185 9741 8219 9775
rect 8253 9741 8287 9775
rect 8321 9741 8355 9775
rect 8389 9741 8423 9775
rect 8457 9741 8491 9775
rect 8525 9741 8559 9775
rect 8593 9741 8627 9775
rect 8661 9741 8695 9775
rect 8729 9741 8763 9775
rect 8797 9741 8831 9775
rect 8865 9741 8899 9775
rect 8933 9741 8967 9775
rect 9001 9741 9035 9775
rect 9069 9741 9103 9775
rect 9137 9741 9171 9775
rect 9205 9741 9239 9775
rect 9273 9741 9307 9775
rect 9341 9741 9375 9775
rect 9409 9741 9443 9775
rect 9477 9741 9511 9775
rect 9545 9741 9579 9775
rect 9613 9741 9647 9775
rect 9681 9741 9715 9775
rect 9749 9741 9783 9775
rect 9817 9741 9851 9775
rect 9885 9741 9919 9775
rect 9953 9741 9987 9775
rect 10021 9741 10055 9775
rect 10089 9741 10123 9775
rect 10157 9741 10191 9775
rect 10225 9741 10259 9775
rect 10293 9741 10327 9775
rect 10361 9741 10395 9775
rect 10429 9741 10463 9775
rect 10497 9741 10531 9775
rect 10565 9741 10599 9775
rect 10633 9741 10667 9775
rect 10701 9741 10735 9775
rect 10769 9741 10803 9775
rect 10837 9741 10871 9775
rect 10905 9741 10939 9775
rect 10973 9741 11007 9775
rect 11041 9741 11075 9775
rect 11109 9741 11143 9775
rect 11177 9741 11211 9775
rect 11245 9741 11279 9775
rect 11313 9741 11347 9775
rect 11381 9741 11415 9775
rect 11449 9741 11483 9775
rect 11517 9741 11551 9775
rect 11585 9741 11619 9775
rect 11653 9741 11687 9775
rect 11721 9741 11755 9775
rect 11789 9741 11823 9775
rect 11857 9741 11891 9775
rect 11925 9741 11959 9775
rect 11993 9741 12027 9775
rect 12061 9741 12095 9775
rect 12129 9741 12163 9775
rect 12197 9741 12231 9775
rect 12265 9741 12299 9775
rect 12333 9741 12367 9775
rect 12401 9741 12435 9775
rect 12469 9741 12503 9775
rect 12537 9741 12571 9775
rect 12605 9741 12639 9775
rect 12673 9741 12707 9775
rect 12741 9741 12775 9775
rect 12809 9741 12843 9775
rect 12877 9741 12911 9775
rect 12945 9741 12979 9775
rect 13013 9741 13047 9775
rect 13081 9741 13115 9775
rect 13149 9741 13183 9775
rect 13217 9741 13251 9775
rect 13285 9741 13319 9775
rect 13353 9741 13387 9775
rect 13421 9741 13455 9775
rect 13489 9741 13523 9775
rect 13557 9741 13591 9775
rect 13625 9741 13659 9775
rect 13693 9741 13727 9775
rect 13761 9741 13795 9775
rect 13829 9741 13863 9775
rect 13897 9741 13931 9775
rect 13965 9741 13999 9775
rect 14033 9741 14067 9775
rect 14101 9741 14135 9775
rect 14169 9741 14203 9775
<< locali >>
rect 245 36534 14724 36574
rect 245 36500 320 36534
rect 354 36533 14724 36534
rect 354 36500 14614 36533
rect 245 36499 14614 36500
rect 14648 36499 14724 36533
rect 245 36465 492 36499
rect 526 36498 560 36499
rect 526 36465 556 36498
rect 594 36465 628 36499
rect 662 36465 696 36499
rect 730 36498 764 36499
rect 798 36498 832 36499
rect 866 36498 900 36499
rect 934 36498 968 36499
rect 1002 36498 1036 36499
rect 1070 36498 1104 36499
rect 1138 36498 1172 36499
rect 1206 36498 1240 36499
rect 734 36465 764 36498
rect 806 36465 832 36498
rect 878 36465 900 36498
rect 950 36465 968 36498
rect 1022 36465 1036 36498
rect 1094 36465 1104 36498
rect 1166 36465 1172 36498
rect 1238 36465 1240 36498
rect 1274 36498 1308 36499
rect 1342 36498 1376 36499
rect 1410 36498 1444 36499
rect 1478 36498 1512 36499
rect 1546 36498 1580 36499
rect 1614 36498 1648 36499
rect 1682 36498 1716 36499
rect 1750 36498 1784 36499
rect 1274 36465 1276 36498
rect 1342 36465 1348 36498
rect 1410 36465 1420 36498
rect 1478 36465 1492 36498
rect 1546 36465 1564 36498
rect 1614 36465 1636 36498
rect 1682 36465 1708 36498
rect 1750 36465 1780 36498
rect 1818 36465 1852 36499
rect 1886 36465 1920 36499
rect 1954 36498 1988 36499
rect 2022 36498 2056 36499
rect 2090 36498 2124 36499
rect 2158 36498 2192 36499
rect 2226 36498 2260 36499
rect 2294 36498 2328 36499
rect 2362 36498 2396 36499
rect 2430 36498 2464 36499
rect 1958 36465 1988 36498
rect 2030 36465 2056 36498
rect 2102 36465 2124 36498
rect 2174 36465 2192 36498
rect 2246 36465 2260 36498
rect 2318 36465 2328 36498
rect 2390 36465 2396 36498
rect 2462 36465 2464 36498
rect 2498 36498 2532 36499
rect 2566 36498 2600 36499
rect 2634 36498 2668 36499
rect 2702 36498 2736 36499
rect 2770 36498 2804 36499
rect 2838 36498 2872 36499
rect 2906 36498 2940 36499
rect 2974 36498 3008 36499
rect 2498 36465 2500 36498
rect 2566 36465 2572 36498
rect 2634 36465 2644 36498
rect 2702 36465 2716 36498
rect 2770 36465 2788 36498
rect 2838 36465 2860 36498
rect 2906 36465 2932 36498
rect 2974 36465 3004 36498
rect 3042 36465 3076 36499
rect 3110 36465 3144 36499
rect 3178 36498 3212 36499
rect 3246 36498 3280 36499
rect 3314 36498 3348 36499
rect 3382 36498 3416 36499
rect 3450 36498 3484 36499
rect 3518 36498 3552 36499
rect 3586 36498 3620 36499
rect 3654 36498 3688 36499
rect 3182 36465 3212 36498
rect 3254 36465 3280 36498
rect 3326 36465 3348 36498
rect 3398 36465 3416 36498
rect 3470 36465 3484 36498
rect 3542 36465 3552 36498
rect 3614 36465 3620 36498
rect 3686 36465 3688 36498
rect 3722 36498 3756 36499
rect 3790 36498 3824 36499
rect 3858 36498 3892 36499
rect 3926 36498 3960 36499
rect 3994 36498 4028 36499
rect 4062 36498 4096 36499
rect 4130 36498 4164 36499
rect 4198 36498 4232 36499
rect 3722 36465 3724 36498
rect 3790 36465 3796 36498
rect 3858 36465 3868 36498
rect 3926 36465 3940 36498
rect 3994 36465 4012 36498
rect 4062 36465 4084 36498
rect 4130 36465 4156 36498
rect 4198 36465 4228 36498
rect 4266 36465 4300 36499
rect 4334 36465 4368 36499
rect 4402 36498 4436 36499
rect 4470 36498 4504 36499
rect 4538 36498 4572 36499
rect 4606 36498 4640 36499
rect 4674 36498 4708 36499
rect 4742 36498 4776 36499
rect 4810 36498 4844 36499
rect 4878 36498 4912 36499
rect 4406 36465 4436 36498
rect 4478 36465 4504 36498
rect 4550 36465 4572 36498
rect 4622 36465 4640 36498
rect 4694 36465 4708 36498
rect 4766 36465 4776 36498
rect 4838 36465 4844 36498
rect 4910 36465 4912 36498
rect 4946 36498 4980 36499
rect 5014 36498 5048 36499
rect 5082 36498 5116 36499
rect 5150 36498 5184 36499
rect 5218 36498 5252 36499
rect 5286 36498 5320 36499
rect 5354 36498 5388 36499
rect 5422 36498 5456 36499
rect 4946 36465 4948 36498
rect 5014 36465 5020 36498
rect 5082 36465 5092 36498
rect 5150 36465 5164 36498
rect 5218 36465 5236 36498
rect 5286 36465 5308 36498
rect 5354 36465 5380 36498
rect 5422 36465 5452 36498
rect 5490 36465 5524 36499
rect 5558 36465 5592 36499
rect 5626 36498 5660 36499
rect 5694 36498 5728 36499
rect 5762 36498 5796 36499
rect 5830 36498 5864 36499
rect 5898 36498 5932 36499
rect 5966 36498 6000 36499
rect 6034 36498 6068 36499
rect 6102 36498 6136 36499
rect 5630 36465 5660 36498
rect 5702 36465 5728 36498
rect 5774 36465 5796 36498
rect 5846 36465 5864 36498
rect 5918 36465 5932 36498
rect 5990 36465 6000 36498
rect 6062 36465 6068 36498
rect 6134 36465 6136 36498
rect 6170 36498 6204 36499
rect 6238 36498 6272 36499
rect 6306 36498 6340 36499
rect 6374 36498 6408 36499
rect 6442 36498 6476 36499
rect 6510 36498 6544 36499
rect 6578 36498 6612 36499
rect 6646 36498 6680 36499
rect 6170 36465 6172 36498
rect 6238 36465 6244 36498
rect 6306 36465 6316 36498
rect 6374 36465 6388 36498
rect 6442 36465 6460 36498
rect 6510 36465 6532 36498
rect 6578 36465 6604 36498
rect 6646 36465 6676 36498
rect 6714 36465 6748 36499
rect 6782 36465 6816 36499
rect 6850 36498 6884 36499
rect 6918 36498 6952 36499
rect 6986 36498 7020 36499
rect 7054 36498 7088 36499
rect 7122 36498 7156 36499
rect 7190 36498 7224 36499
rect 7258 36498 7292 36499
rect 7326 36498 7360 36499
rect 6854 36465 6884 36498
rect 6926 36465 6952 36498
rect 6998 36465 7020 36498
rect 7070 36465 7088 36498
rect 7142 36465 7156 36498
rect 7214 36465 7224 36498
rect 7286 36465 7292 36498
rect 7358 36465 7360 36498
rect 7394 36498 7428 36499
rect 7462 36498 7496 36499
rect 7530 36498 7564 36499
rect 7598 36498 7632 36499
rect 7666 36498 7700 36499
rect 7734 36498 7768 36499
rect 7802 36498 7836 36499
rect 7870 36498 7904 36499
rect 7394 36465 7396 36498
rect 7462 36465 7468 36498
rect 7530 36465 7540 36498
rect 7598 36465 7612 36498
rect 7666 36465 7684 36498
rect 7734 36465 7756 36498
rect 7802 36465 7828 36498
rect 7870 36465 7900 36498
rect 7938 36465 7972 36499
rect 8006 36465 8040 36499
rect 8074 36498 8108 36499
rect 8142 36498 8176 36499
rect 8210 36498 8244 36499
rect 8278 36498 8312 36499
rect 8346 36498 8380 36499
rect 8414 36498 8448 36499
rect 8482 36498 8516 36499
rect 8550 36498 8584 36499
rect 8078 36465 8108 36498
rect 8150 36465 8176 36498
rect 8222 36465 8244 36498
rect 8294 36465 8312 36498
rect 8366 36465 8380 36498
rect 8438 36465 8448 36498
rect 8510 36465 8516 36498
rect 8582 36465 8584 36498
rect 8618 36498 8652 36499
rect 8686 36498 8720 36499
rect 8754 36498 8788 36499
rect 8822 36498 8856 36499
rect 8890 36498 8924 36499
rect 8958 36498 8992 36499
rect 9026 36498 9060 36499
rect 9094 36498 9128 36499
rect 8618 36465 8620 36498
rect 8686 36465 8692 36498
rect 8754 36465 8764 36498
rect 8822 36465 8836 36498
rect 8890 36465 8908 36498
rect 8958 36465 8980 36498
rect 9026 36465 9052 36498
rect 9094 36465 9124 36498
rect 9162 36465 9196 36499
rect 9230 36465 9264 36499
rect 9298 36498 9332 36499
rect 9366 36498 9400 36499
rect 9434 36498 9468 36499
rect 9502 36498 9536 36499
rect 9570 36498 9604 36499
rect 9638 36498 9672 36499
rect 9706 36498 9740 36499
rect 9774 36498 9808 36499
rect 9302 36465 9332 36498
rect 9374 36465 9400 36498
rect 9446 36465 9468 36498
rect 9518 36465 9536 36498
rect 9590 36465 9604 36498
rect 9662 36465 9672 36498
rect 9734 36465 9740 36498
rect 9806 36465 9808 36498
rect 9842 36498 9876 36499
rect 9910 36498 9944 36499
rect 9978 36498 10012 36499
rect 10046 36498 10080 36499
rect 10114 36498 10148 36499
rect 10182 36498 10216 36499
rect 10250 36498 10284 36499
rect 10318 36498 10352 36499
rect 9842 36465 9844 36498
rect 9910 36465 9916 36498
rect 9978 36465 9988 36498
rect 10046 36465 10060 36498
rect 10114 36465 10132 36498
rect 10182 36465 10204 36498
rect 10250 36465 10276 36498
rect 10318 36465 10348 36498
rect 10386 36465 10420 36499
rect 10454 36465 10488 36499
rect 10522 36498 10556 36499
rect 10590 36498 10624 36499
rect 10658 36498 10692 36499
rect 10726 36498 10760 36499
rect 10794 36498 10828 36499
rect 10862 36498 10896 36499
rect 10930 36498 10964 36499
rect 10998 36498 11032 36499
rect 10526 36465 10556 36498
rect 10598 36465 10624 36498
rect 10670 36465 10692 36498
rect 10742 36465 10760 36498
rect 10814 36465 10828 36498
rect 10886 36465 10896 36498
rect 10958 36465 10964 36498
rect 11030 36465 11032 36498
rect 11066 36498 11100 36499
rect 11134 36498 11168 36499
rect 11202 36498 11236 36499
rect 11270 36498 11304 36499
rect 11338 36498 11372 36499
rect 11406 36498 11440 36499
rect 11474 36498 11508 36499
rect 11542 36498 11576 36499
rect 11066 36465 11068 36498
rect 11134 36465 11140 36498
rect 11202 36465 11212 36498
rect 11270 36465 11284 36498
rect 11338 36465 11356 36498
rect 11406 36465 11428 36498
rect 11474 36465 11500 36498
rect 11542 36465 11572 36498
rect 11610 36465 11644 36499
rect 11678 36465 11712 36499
rect 11746 36498 11780 36499
rect 11814 36498 11848 36499
rect 11882 36498 11916 36499
rect 11950 36498 11984 36499
rect 12018 36498 12052 36499
rect 12086 36498 12120 36499
rect 12154 36498 12188 36499
rect 12222 36498 12256 36499
rect 11750 36465 11780 36498
rect 11822 36465 11848 36498
rect 11894 36465 11916 36498
rect 11966 36465 11984 36498
rect 12038 36465 12052 36498
rect 12110 36465 12120 36498
rect 12182 36465 12188 36498
rect 12254 36465 12256 36498
rect 12290 36498 12324 36499
rect 12358 36498 12392 36499
rect 12426 36498 12460 36499
rect 12494 36498 12528 36499
rect 12562 36498 12596 36499
rect 12630 36498 12664 36499
rect 12698 36498 12732 36499
rect 12766 36498 12800 36499
rect 12290 36465 12292 36498
rect 12358 36465 12364 36498
rect 12426 36465 12436 36498
rect 12494 36465 12508 36498
rect 12562 36465 12580 36498
rect 12630 36465 12652 36498
rect 12698 36465 12724 36498
rect 12766 36465 12796 36498
rect 12834 36465 12868 36499
rect 12902 36465 12936 36499
rect 12970 36498 13004 36499
rect 13038 36498 13072 36499
rect 13106 36498 13140 36499
rect 13174 36498 13208 36499
rect 13242 36498 13276 36499
rect 13310 36498 13344 36499
rect 13378 36498 13412 36499
rect 13446 36498 13480 36499
rect 12974 36465 13004 36498
rect 13046 36465 13072 36498
rect 13118 36465 13140 36498
rect 13190 36465 13208 36498
rect 13262 36465 13276 36498
rect 13334 36465 13344 36498
rect 13406 36465 13412 36498
rect 13478 36465 13480 36498
rect 13514 36498 13548 36499
rect 13582 36498 13616 36499
rect 13650 36498 13684 36499
rect 13718 36498 13752 36499
rect 13786 36498 13820 36499
rect 13854 36498 13888 36499
rect 13922 36498 13956 36499
rect 13990 36498 14024 36499
rect 13514 36465 13516 36498
rect 13582 36465 13588 36498
rect 13650 36465 13660 36498
rect 13718 36465 13732 36498
rect 13786 36465 13804 36498
rect 13854 36465 13876 36498
rect 13922 36465 13948 36498
rect 13990 36465 14020 36498
rect 14058 36465 14092 36499
rect 14126 36465 14160 36499
rect 14194 36498 14228 36499
rect 14262 36498 14296 36499
rect 14330 36498 14364 36499
rect 14398 36498 14432 36499
rect 14198 36465 14228 36498
rect 14270 36465 14296 36498
rect 14342 36465 14364 36498
rect 14414 36465 14432 36498
rect 14466 36465 14724 36499
rect 245 36464 556 36465
rect 590 36464 628 36465
rect 662 36464 700 36465
rect 734 36464 772 36465
rect 806 36464 844 36465
rect 878 36464 916 36465
rect 950 36464 988 36465
rect 1022 36464 1060 36465
rect 1094 36464 1132 36465
rect 1166 36464 1204 36465
rect 1238 36464 1276 36465
rect 1310 36464 1348 36465
rect 1382 36464 1420 36465
rect 1454 36464 1492 36465
rect 1526 36464 1564 36465
rect 1598 36464 1636 36465
rect 1670 36464 1708 36465
rect 1742 36464 1780 36465
rect 1814 36464 1852 36465
rect 1886 36464 1924 36465
rect 1958 36464 1996 36465
rect 2030 36464 2068 36465
rect 2102 36464 2140 36465
rect 2174 36464 2212 36465
rect 2246 36464 2284 36465
rect 2318 36464 2356 36465
rect 2390 36464 2428 36465
rect 2462 36464 2500 36465
rect 2534 36464 2572 36465
rect 2606 36464 2644 36465
rect 2678 36464 2716 36465
rect 2750 36464 2788 36465
rect 2822 36464 2860 36465
rect 2894 36464 2932 36465
rect 2966 36464 3004 36465
rect 3038 36464 3076 36465
rect 3110 36464 3148 36465
rect 3182 36464 3220 36465
rect 3254 36464 3292 36465
rect 3326 36464 3364 36465
rect 3398 36464 3436 36465
rect 3470 36464 3508 36465
rect 3542 36464 3580 36465
rect 3614 36464 3652 36465
rect 3686 36464 3724 36465
rect 3758 36464 3796 36465
rect 3830 36464 3868 36465
rect 3902 36464 3940 36465
rect 3974 36464 4012 36465
rect 4046 36464 4084 36465
rect 4118 36464 4156 36465
rect 4190 36464 4228 36465
rect 4262 36464 4300 36465
rect 4334 36464 4372 36465
rect 4406 36464 4444 36465
rect 4478 36464 4516 36465
rect 4550 36464 4588 36465
rect 4622 36464 4660 36465
rect 4694 36464 4732 36465
rect 4766 36464 4804 36465
rect 4838 36464 4876 36465
rect 4910 36464 4948 36465
rect 4982 36464 5020 36465
rect 5054 36464 5092 36465
rect 5126 36464 5164 36465
rect 5198 36464 5236 36465
rect 5270 36464 5308 36465
rect 5342 36464 5380 36465
rect 5414 36464 5452 36465
rect 5486 36464 5524 36465
rect 5558 36464 5596 36465
rect 5630 36464 5668 36465
rect 5702 36464 5740 36465
rect 5774 36464 5812 36465
rect 5846 36464 5884 36465
rect 5918 36464 5956 36465
rect 5990 36464 6028 36465
rect 6062 36464 6100 36465
rect 6134 36464 6172 36465
rect 6206 36464 6244 36465
rect 6278 36464 6316 36465
rect 6350 36464 6388 36465
rect 6422 36464 6460 36465
rect 6494 36464 6532 36465
rect 6566 36464 6604 36465
rect 6638 36464 6676 36465
rect 6710 36464 6748 36465
rect 6782 36464 6820 36465
rect 6854 36464 6892 36465
rect 6926 36464 6964 36465
rect 6998 36464 7036 36465
rect 7070 36464 7108 36465
rect 7142 36464 7180 36465
rect 7214 36464 7252 36465
rect 7286 36464 7324 36465
rect 7358 36464 7396 36465
rect 7430 36464 7468 36465
rect 7502 36464 7540 36465
rect 7574 36464 7612 36465
rect 7646 36464 7684 36465
rect 7718 36464 7756 36465
rect 7790 36464 7828 36465
rect 7862 36464 7900 36465
rect 7934 36464 7972 36465
rect 8006 36464 8044 36465
rect 8078 36464 8116 36465
rect 8150 36464 8188 36465
rect 8222 36464 8260 36465
rect 8294 36464 8332 36465
rect 8366 36464 8404 36465
rect 8438 36464 8476 36465
rect 8510 36464 8548 36465
rect 8582 36464 8620 36465
rect 8654 36464 8692 36465
rect 8726 36464 8764 36465
rect 8798 36464 8836 36465
rect 8870 36464 8908 36465
rect 8942 36464 8980 36465
rect 9014 36464 9052 36465
rect 9086 36464 9124 36465
rect 9158 36464 9196 36465
rect 9230 36464 9268 36465
rect 9302 36464 9340 36465
rect 9374 36464 9412 36465
rect 9446 36464 9484 36465
rect 9518 36464 9556 36465
rect 9590 36464 9628 36465
rect 9662 36464 9700 36465
rect 9734 36464 9772 36465
rect 9806 36464 9844 36465
rect 9878 36464 9916 36465
rect 9950 36464 9988 36465
rect 10022 36464 10060 36465
rect 10094 36464 10132 36465
rect 10166 36464 10204 36465
rect 10238 36464 10276 36465
rect 10310 36464 10348 36465
rect 10382 36464 10420 36465
rect 10454 36464 10492 36465
rect 10526 36464 10564 36465
rect 10598 36464 10636 36465
rect 10670 36464 10708 36465
rect 10742 36464 10780 36465
rect 10814 36464 10852 36465
rect 10886 36464 10924 36465
rect 10958 36464 10996 36465
rect 11030 36464 11068 36465
rect 11102 36464 11140 36465
rect 11174 36464 11212 36465
rect 11246 36464 11284 36465
rect 11318 36464 11356 36465
rect 11390 36464 11428 36465
rect 11462 36464 11500 36465
rect 11534 36464 11572 36465
rect 11606 36464 11644 36465
rect 11678 36464 11716 36465
rect 11750 36464 11788 36465
rect 11822 36464 11860 36465
rect 11894 36464 11932 36465
rect 11966 36464 12004 36465
rect 12038 36464 12076 36465
rect 12110 36464 12148 36465
rect 12182 36464 12220 36465
rect 12254 36464 12292 36465
rect 12326 36464 12364 36465
rect 12398 36464 12436 36465
rect 12470 36464 12508 36465
rect 12542 36464 12580 36465
rect 12614 36464 12652 36465
rect 12686 36464 12724 36465
rect 12758 36464 12796 36465
rect 12830 36464 12868 36465
rect 12902 36464 12940 36465
rect 12974 36464 13012 36465
rect 13046 36464 13084 36465
rect 13118 36464 13156 36465
rect 13190 36464 13228 36465
rect 13262 36464 13300 36465
rect 13334 36464 13372 36465
rect 13406 36464 13444 36465
rect 13478 36464 13516 36465
rect 13550 36464 13588 36465
rect 13622 36464 13660 36465
rect 13694 36464 13732 36465
rect 13766 36464 13804 36465
rect 13838 36464 13876 36465
rect 13910 36464 13948 36465
rect 13982 36464 14020 36465
rect 14054 36464 14092 36465
rect 14126 36464 14164 36465
rect 14198 36464 14236 36465
rect 14270 36464 14308 36465
rect 14342 36464 14380 36465
rect 14414 36464 14724 36465
rect 245 36462 14724 36464
rect 245 36428 320 36462
rect 354 36461 14724 36462
rect 354 36428 14614 36461
rect 245 36427 14614 36428
rect 14648 36427 14724 36461
rect 245 36389 14724 36427
rect 245 36335 430 36389
rect 245 36301 322 36335
rect 356 36301 430 36335
rect 245 36267 430 36301
rect 245 36265 322 36267
rect 245 36231 320 36265
rect 356 36233 430 36267
rect 354 36231 430 36233
rect 245 36199 430 36231
rect 14539 36327 14724 36389
rect 14539 36293 14609 36327
rect 14643 36293 14724 36327
rect 14539 36262 14724 36293
rect 14539 36259 14614 36262
rect 14539 36225 14609 36259
rect 14648 36228 14724 36262
rect 14643 36225 14724 36228
rect 245 36193 322 36199
rect 245 36159 320 36193
rect 356 36165 430 36199
rect 354 36159 430 36165
rect 245 36131 430 36159
rect 245 36121 322 36131
rect 245 36087 320 36121
rect 356 36097 430 36131
rect 354 36087 430 36097
rect 245 36063 430 36087
rect 245 36049 322 36063
rect 245 36015 320 36049
rect 356 36029 430 36063
rect 354 36015 430 36029
rect 245 35995 430 36015
rect 245 35977 322 35995
rect 245 35943 320 35977
rect 356 35961 430 35995
rect 354 35943 430 35961
rect 245 35927 430 35943
rect 245 35905 322 35927
rect 245 35871 320 35905
rect 356 35893 430 35927
rect 354 35871 430 35893
rect 245 35859 430 35871
rect 245 35833 322 35859
rect 245 35799 320 35833
rect 356 35825 430 35859
rect 354 35799 430 35825
rect 245 35791 430 35799
rect 245 35761 322 35791
rect 245 35727 320 35761
rect 356 35757 430 35791
rect 354 35727 430 35757
rect 245 35723 430 35727
rect 245 35689 322 35723
rect 356 35689 430 35723
rect 245 35655 320 35689
rect 354 35655 430 35689
rect 245 35621 322 35655
rect 356 35621 430 35655
rect 245 35617 430 35621
rect 245 35583 320 35617
rect 354 35587 430 35617
rect 245 35553 322 35583
rect 356 35553 430 35587
rect 245 35545 430 35553
rect 245 35511 320 35545
rect 354 35519 430 35545
rect 245 35485 322 35511
rect 356 35485 430 35519
rect 245 35473 430 35485
rect 245 35439 320 35473
rect 354 35451 430 35473
rect 245 35417 322 35439
rect 356 35417 430 35451
rect 245 35401 430 35417
rect 245 35367 320 35401
rect 354 35383 430 35401
rect 245 35349 322 35367
rect 356 35349 430 35383
rect 245 35329 430 35349
rect 245 35295 320 35329
rect 354 35315 430 35329
rect 245 35281 322 35295
rect 356 35281 430 35315
rect 245 35257 430 35281
rect 245 35223 320 35257
rect 354 35247 430 35257
rect 245 35213 322 35223
rect 356 35213 430 35247
rect 245 35185 430 35213
rect 245 35151 320 35185
rect 354 35179 430 35185
rect 245 35145 322 35151
rect 356 35145 430 35179
rect 245 35113 430 35145
rect 245 35079 320 35113
rect 354 35111 430 35113
rect 245 35077 322 35079
rect 356 35077 430 35111
rect 245 35043 430 35077
rect 245 35041 322 35043
rect 245 35007 320 35041
rect 356 35009 430 35043
rect 354 35007 430 35009
rect 245 34975 430 35007
rect 245 34969 322 34975
rect 245 34935 320 34969
rect 356 34941 430 34975
rect 354 34935 430 34941
rect 245 34907 430 34935
rect 245 34897 322 34907
rect 245 34863 320 34897
rect 356 34873 430 34907
rect 354 34863 430 34873
rect 245 34839 430 34863
rect 245 34825 322 34839
rect 245 34791 320 34825
rect 356 34805 430 34839
rect 354 34791 430 34805
rect 245 34771 430 34791
rect 245 34753 322 34771
rect 245 34719 320 34753
rect 356 34737 430 34771
rect 354 34719 430 34737
rect 245 34703 430 34719
rect 245 34681 322 34703
rect 245 34647 320 34681
rect 356 34669 430 34703
rect 354 34647 430 34669
rect 245 34635 430 34647
rect 245 34609 322 34635
rect 245 34575 320 34609
rect 356 34601 430 34635
rect 354 34575 430 34601
rect 245 34567 430 34575
rect 245 34537 322 34567
rect 245 34503 320 34537
rect 356 34533 430 34567
rect 354 34503 430 34533
rect 245 34499 430 34503
rect 245 34465 322 34499
rect 356 34465 430 34499
rect 245 34431 320 34465
rect 354 34431 430 34465
rect 245 34397 322 34431
rect 356 34397 430 34431
rect 245 34393 430 34397
rect 245 34359 320 34393
rect 354 34363 430 34393
rect 245 34329 322 34359
rect 356 34329 430 34363
rect 245 34321 430 34329
rect 245 34287 320 34321
rect 354 34295 430 34321
rect 245 34261 322 34287
rect 356 34261 430 34295
rect 245 34249 430 34261
rect 245 34215 320 34249
rect 354 34227 430 34249
rect 245 34193 322 34215
rect 356 34193 430 34227
rect 245 34177 430 34193
rect 245 34143 320 34177
rect 354 34159 430 34177
rect 245 34125 322 34143
rect 356 34125 430 34159
rect 245 34105 430 34125
rect 245 34071 320 34105
rect 354 34091 430 34105
rect 245 34057 322 34071
rect 356 34057 430 34091
rect 245 34033 430 34057
rect 245 33999 320 34033
rect 354 34023 430 34033
rect 245 33989 322 33999
rect 356 33989 430 34023
rect 245 33961 430 33989
rect 245 33927 320 33961
rect 354 33955 430 33961
rect 245 33921 322 33927
rect 356 33921 430 33955
rect 245 33889 430 33921
rect 245 33855 320 33889
rect 354 33887 430 33889
rect 245 33853 322 33855
rect 356 33853 430 33887
rect 245 33819 430 33853
rect 245 33817 322 33819
rect 245 33783 320 33817
rect 356 33785 430 33819
rect 354 33783 430 33785
rect 245 33751 430 33783
rect 245 33745 322 33751
rect 245 33711 320 33745
rect 356 33717 430 33751
rect 354 33711 430 33717
rect 245 33683 430 33711
rect 245 33673 322 33683
rect 245 33639 320 33673
rect 356 33649 430 33683
rect 354 33639 430 33649
rect 245 33615 430 33639
rect 245 33601 322 33615
rect 245 33567 320 33601
rect 356 33581 430 33615
rect 354 33567 430 33581
rect 245 33547 430 33567
rect 245 33529 322 33547
rect 245 33495 320 33529
rect 356 33513 430 33547
rect 354 33495 430 33513
rect 245 33479 430 33495
rect 245 33457 322 33479
rect 245 33423 320 33457
rect 356 33445 430 33479
rect 354 33423 430 33445
rect 245 33411 430 33423
rect 245 33385 322 33411
rect 245 33351 320 33385
rect 356 33377 430 33411
rect 354 33351 430 33377
rect 245 33343 430 33351
rect 245 33313 322 33343
rect 245 33279 320 33313
rect 356 33309 430 33343
rect 354 33279 430 33309
rect 245 33275 430 33279
rect 245 33241 322 33275
rect 356 33241 430 33275
rect 245 33207 320 33241
rect 354 33207 430 33241
rect 245 33173 322 33207
rect 356 33173 430 33207
rect 245 33169 430 33173
rect 245 33135 320 33169
rect 354 33139 430 33169
rect 245 33105 322 33135
rect 356 33105 430 33139
rect 245 33097 430 33105
rect 245 33063 320 33097
rect 354 33071 430 33097
rect 245 33037 322 33063
rect 356 33037 430 33071
rect 245 33025 430 33037
rect 245 32991 320 33025
rect 354 33003 430 33025
rect 245 32969 322 32991
rect 356 32969 430 33003
rect 245 32953 430 32969
rect 245 32919 320 32953
rect 354 32935 430 32953
rect 245 32901 322 32919
rect 356 32901 430 32935
rect 245 32881 430 32901
rect 245 32847 320 32881
rect 354 32867 430 32881
rect 245 32833 322 32847
rect 356 32833 430 32867
rect 245 32809 430 32833
rect 245 32775 320 32809
rect 354 32799 430 32809
rect 245 32765 322 32775
rect 356 32765 430 32799
rect 245 32737 430 32765
rect 245 32703 320 32737
rect 354 32731 430 32737
rect 245 32697 322 32703
rect 356 32697 430 32731
rect 245 32665 430 32697
rect 245 32631 320 32665
rect 354 32663 430 32665
rect 245 32629 322 32631
rect 356 32629 430 32663
rect 245 32595 430 32629
rect 245 32593 322 32595
rect 245 32559 320 32593
rect 356 32561 430 32595
rect 354 32559 430 32561
rect 245 32527 430 32559
rect 245 32521 322 32527
rect 245 32487 320 32521
rect 356 32493 430 32527
rect 354 32487 430 32493
rect 245 32459 430 32487
rect 245 32449 322 32459
rect 245 32415 320 32449
rect 356 32425 430 32459
rect 354 32415 430 32425
rect 245 32391 430 32415
rect 245 32377 322 32391
rect 245 32343 320 32377
rect 356 32357 430 32391
rect 354 32343 430 32357
rect 245 32323 430 32343
rect 245 32305 322 32323
rect 245 32271 320 32305
rect 356 32289 430 32323
rect 354 32271 430 32289
rect 245 32255 430 32271
rect 245 32233 322 32255
rect 245 32199 320 32233
rect 356 32221 430 32255
rect 354 32199 430 32221
rect 245 32187 430 32199
rect 245 32161 322 32187
rect 245 32127 320 32161
rect 356 32153 430 32187
rect 354 32127 430 32153
rect 245 32119 430 32127
rect 245 32089 322 32119
rect 245 32055 320 32089
rect 356 32085 430 32119
rect 354 32055 430 32085
rect 245 32051 430 32055
rect 245 32017 322 32051
rect 356 32017 430 32051
rect 245 31983 320 32017
rect 354 31983 430 32017
rect 245 31949 322 31983
rect 356 31949 430 31983
rect 245 31945 430 31949
rect 245 31911 320 31945
rect 354 31915 430 31945
rect 245 31881 322 31911
rect 356 31881 430 31915
rect 245 31873 430 31881
rect 245 31839 320 31873
rect 354 31847 430 31873
rect 245 31813 322 31839
rect 356 31813 430 31847
rect 245 31801 430 31813
rect 245 31767 320 31801
rect 354 31779 430 31801
rect 245 31745 322 31767
rect 356 31745 430 31779
rect 245 31729 430 31745
rect 245 31695 320 31729
rect 354 31711 430 31729
rect 245 31677 322 31695
rect 356 31677 430 31711
rect 245 31657 430 31677
rect 245 31623 320 31657
rect 354 31643 430 31657
rect 245 31609 322 31623
rect 356 31609 430 31643
rect 245 31585 430 31609
rect 245 31551 320 31585
rect 354 31575 430 31585
rect 245 31541 322 31551
rect 356 31541 430 31575
rect 245 31513 430 31541
rect 245 31479 320 31513
rect 354 31507 430 31513
rect 245 31473 322 31479
rect 356 31473 430 31507
rect 245 31441 430 31473
rect 245 31407 320 31441
rect 354 31439 430 31441
rect 245 31405 322 31407
rect 356 31405 430 31439
rect 245 31371 430 31405
rect 245 31369 322 31371
rect 245 31335 320 31369
rect 356 31337 430 31371
rect 354 31335 430 31337
rect 245 31303 430 31335
rect 245 31297 322 31303
rect 245 31263 320 31297
rect 356 31269 430 31303
rect 354 31263 430 31269
rect 245 31235 430 31263
rect 245 31225 322 31235
rect 245 31191 320 31225
rect 356 31201 430 31235
rect 354 31191 430 31201
rect 245 31167 430 31191
rect 245 31153 322 31167
rect 245 31119 320 31153
rect 356 31133 430 31167
rect 354 31119 430 31133
rect 245 31099 430 31119
rect 245 31081 322 31099
rect 245 31047 320 31081
rect 356 31065 430 31099
rect 354 31047 430 31065
rect 245 31031 430 31047
rect 245 31009 322 31031
rect 245 30975 320 31009
rect 356 30997 430 31031
rect 354 30975 430 30997
rect 245 30963 430 30975
rect 245 30937 322 30963
rect 245 30903 320 30937
rect 356 30929 430 30963
rect 354 30903 430 30929
rect 245 30895 430 30903
rect 245 30865 322 30895
rect 245 30831 320 30865
rect 356 30861 430 30895
rect 354 30831 430 30861
rect 245 30827 430 30831
rect 245 30793 322 30827
rect 356 30793 430 30827
rect 245 30759 320 30793
rect 354 30759 430 30793
rect 245 30725 322 30759
rect 356 30725 430 30759
rect 245 30721 430 30725
rect 245 30687 320 30721
rect 354 30691 430 30721
rect 245 30657 322 30687
rect 356 30657 430 30691
rect 245 30649 430 30657
rect 245 30615 320 30649
rect 354 30623 430 30649
rect 245 30589 322 30615
rect 356 30589 430 30623
rect 245 30577 430 30589
rect 245 30543 320 30577
rect 354 30555 430 30577
rect 245 30521 322 30543
rect 356 30521 430 30555
rect 245 30505 430 30521
rect 245 30471 320 30505
rect 354 30487 430 30505
rect 245 30453 322 30471
rect 356 30453 430 30487
rect 245 30433 430 30453
rect 245 30399 320 30433
rect 354 30419 430 30433
rect 245 30385 322 30399
rect 356 30385 430 30419
rect 245 30361 430 30385
rect 245 30327 320 30361
rect 354 30351 430 30361
rect 245 30317 322 30327
rect 356 30317 430 30351
rect 245 30289 430 30317
rect 245 30255 320 30289
rect 354 30283 430 30289
rect 245 30249 322 30255
rect 356 30249 430 30283
rect 245 30217 430 30249
rect 245 30183 320 30217
rect 354 30215 430 30217
rect 245 30181 322 30183
rect 356 30181 430 30215
rect 245 30147 430 30181
rect 245 30145 322 30147
rect 245 30111 320 30145
rect 356 30113 430 30147
rect 354 30111 430 30113
rect 245 30079 430 30111
rect 245 30073 322 30079
rect 245 30039 320 30073
rect 356 30045 430 30079
rect 354 30039 430 30045
rect 245 30011 430 30039
rect 245 30001 322 30011
rect 245 29967 320 30001
rect 356 29977 430 30011
rect 354 29967 430 29977
rect 245 29943 430 29967
rect 245 29929 322 29943
rect 245 29895 320 29929
rect 356 29909 430 29943
rect 354 29895 430 29909
rect 245 29875 430 29895
rect 245 29857 322 29875
rect 245 29823 320 29857
rect 356 29841 430 29875
rect 354 29823 430 29841
rect 245 29807 430 29823
rect 245 29785 322 29807
rect 245 29751 320 29785
rect 356 29773 430 29807
rect 354 29751 430 29773
rect 245 29739 430 29751
rect 245 29713 322 29739
rect 245 29679 320 29713
rect 356 29705 430 29739
rect 354 29679 430 29705
rect 245 29671 430 29679
rect 245 29641 322 29671
rect 245 29607 320 29641
rect 356 29637 430 29671
rect 354 29607 430 29637
rect 245 29603 430 29607
rect 245 29569 322 29603
rect 356 29569 430 29603
rect 245 29535 320 29569
rect 354 29535 430 29569
rect 245 29501 322 29535
rect 356 29501 430 29535
rect 245 29497 430 29501
rect 245 29463 320 29497
rect 354 29467 430 29497
rect 245 29433 322 29463
rect 356 29433 430 29467
rect 245 29425 430 29433
rect 245 29391 320 29425
rect 354 29399 430 29425
rect 245 29365 322 29391
rect 356 29365 430 29399
rect 245 29353 430 29365
rect 245 29319 320 29353
rect 354 29331 430 29353
rect 245 29297 322 29319
rect 356 29297 430 29331
rect 245 29281 430 29297
rect 245 29247 320 29281
rect 354 29263 430 29281
rect 245 29229 322 29247
rect 356 29229 430 29263
rect 245 29209 430 29229
rect 245 29175 320 29209
rect 354 29195 430 29209
rect 245 29161 322 29175
rect 356 29161 430 29195
rect 245 29137 430 29161
rect 245 29103 320 29137
rect 354 29127 430 29137
rect 245 29093 322 29103
rect 356 29093 430 29127
rect 245 29065 430 29093
rect 245 29031 320 29065
rect 354 29059 430 29065
rect 245 29025 322 29031
rect 356 29025 430 29059
rect 245 28993 430 29025
rect 245 28959 320 28993
rect 354 28991 430 28993
rect 245 28957 322 28959
rect 356 28957 430 28991
rect 245 28923 430 28957
rect 245 28921 322 28923
rect 245 28887 320 28921
rect 356 28889 430 28923
rect 354 28887 430 28889
rect 245 28855 430 28887
rect 245 28849 322 28855
rect 245 28815 320 28849
rect 356 28821 430 28855
rect 354 28815 430 28821
rect 245 28787 430 28815
rect 245 28777 322 28787
rect 245 28743 320 28777
rect 356 28753 430 28787
rect 354 28743 430 28753
rect 245 28719 430 28743
rect 245 28705 322 28719
rect 245 28671 320 28705
rect 356 28685 430 28719
rect 354 28671 430 28685
rect 245 28651 430 28671
rect 245 28633 322 28651
rect 245 28599 320 28633
rect 356 28617 430 28651
rect 354 28599 430 28617
rect 245 28583 430 28599
rect 245 28561 322 28583
rect 245 28527 320 28561
rect 356 28549 430 28583
rect 354 28527 430 28549
rect 245 28515 430 28527
rect 245 28489 322 28515
rect 245 28455 320 28489
rect 356 28481 430 28515
rect 354 28455 430 28481
rect 245 28447 430 28455
rect 245 28417 322 28447
rect 245 28383 320 28417
rect 356 28413 430 28447
rect 354 28383 430 28413
rect 245 28379 430 28383
rect 245 28345 322 28379
rect 356 28345 430 28379
rect 245 28311 320 28345
rect 354 28311 430 28345
rect 245 28277 322 28311
rect 356 28277 430 28311
rect 245 28273 430 28277
rect 245 28239 320 28273
rect 354 28243 430 28273
rect 245 28209 322 28239
rect 356 28209 430 28243
rect 245 28201 430 28209
rect 245 28167 320 28201
rect 354 28175 430 28201
rect 245 28141 322 28167
rect 356 28141 430 28175
rect 245 28129 430 28141
rect 245 28095 320 28129
rect 354 28107 430 28129
rect 245 28073 322 28095
rect 356 28073 430 28107
rect 245 28057 430 28073
rect 245 28023 320 28057
rect 354 28039 430 28057
rect 245 28005 322 28023
rect 356 28005 430 28039
rect 245 27985 430 28005
rect 245 27951 320 27985
rect 354 27971 430 27985
rect 245 27937 322 27951
rect 356 27937 430 27971
rect 245 27913 430 27937
rect 245 27879 320 27913
rect 354 27903 430 27913
rect 245 27869 322 27879
rect 356 27869 430 27903
rect 245 27841 430 27869
rect 245 27807 320 27841
rect 354 27835 430 27841
rect 245 27801 322 27807
rect 356 27801 430 27835
rect 245 27769 430 27801
rect 245 27735 320 27769
rect 354 27767 430 27769
rect 245 27733 322 27735
rect 356 27733 430 27767
rect 245 27699 430 27733
rect 245 27697 322 27699
rect 245 27663 320 27697
rect 356 27665 430 27699
rect 354 27663 430 27665
rect 245 27631 430 27663
rect 245 27625 322 27631
rect 245 27591 320 27625
rect 356 27597 430 27631
rect 354 27591 430 27597
rect 245 27563 430 27591
rect 245 27553 322 27563
rect 245 27519 320 27553
rect 356 27529 430 27563
rect 354 27519 430 27529
rect 245 27495 430 27519
rect 245 27481 322 27495
rect 245 27447 320 27481
rect 356 27461 430 27495
rect 354 27447 430 27461
rect 245 27427 430 27447
rect 245 27409 322 27427
rect 245 27375 320 27409
rect 356 27393 430 27427
rect 354 27375 430 27393
rect 245 27359 430 27375
rect 245 27337 322 27359
rect 245 27303 320 27337
rect 356 27325 430 27359
rect 354 27303 430 27325
rect 245 27291 430 27303
rect 245 27265 322 27291
rect 245 27231 320 27265
rect 356 27257 430 27291
rect 354 27231 430 27257
rect 245 27223 430 27231
rect 245 27193 322 27223
rect 245 27159 320 27193
rect 356 27189 430 27223
rect 354 27159 430 27189
rect 245 27155 430 27159
rect 245 27121 322 27155
rect 356 27121 430 27155
rect 245 27087 320 27121
rect 354 27087 430 27121
rect 245 27053 322 27087
rect 356 27053 430 27087
rect 245 27049 430 27053
rect 245 27015 320 27049
rect 354 27019 430 27049
rect 245 26985 322 27015
rect 356 26985 430 27019
rect 245 26977 430 26985
rect 245 26943 320 26977
rect 354 26951 430 26977
rect 245 26917 322 26943
rect 356 26917 430 26951
rect 245 26905 430 26917
rect 245 26871 320 26905
rect 354 26883 430 26905
rect 245 26849 322 26871
rect 356 26849 430 26883
rect 245 26833 430 26849
rect 245 26799 320 26833
rect 354 26815 430 26833
rect 245 26781 322 26799
rect 356 26781 430 26815
rect 245 26761 430 26781
rect 245 26727 320 26761
rect 354 26747 430 26761
rect 245 26713 322 26727
rect 356 26713 430 26747
rect 245 26689 430 26713
rect 245 26655 320 26689
rect 354 26679 430 26689
rect 245 26645 322 26655
rect 356 26645 430 26679
rect 245 26617 430 26645
rect 245 26583 320 26617
rect 354 26611 430 26617
rect 245 26577 322 26583
rect 356 26577 430 26611
rect 245 26545 430 26577
rect 245 26511 320 26545
rect 354 26543 430 26545
rect 245 26509 322 26511
rect 356 26509 430 26543
rect 245 26475 430 26509
rect 245 26473 322 26475
rect 245 26439 320 26473
rect 356 26441 430 26475
rect 354 26439 430 26441
rect 245 26407 430 26439
rect 245 26401 322 26407
rect 245 26367 320 26401
rect 356 26373 430 26407
rect 354 26367 430 26373
rect 245 26339 430 26367
rect 245 26329 322 26339
rect 245 26295 320 26329
rect 356 26305 430 26339
rect 354 26295 430 26305
rect 245 26271 430 26295
rect 245 26257 322 26271
rect 245 26223 320 26257
rect 356 26237 430 26271
rect 354 26223 430 26237
rect 245 26203 430 26223
rect 245 26185 322 26203
rect 245 26151 320 26185
rect 356 26169 430 26203
rect 354 26151 430 26169
rect 245 26135 430 26151
rect 245 26113 322 26135
rect 245 26079 320 26113
rect 356 26101 430 26135
rect 354 26079 430 26101
rect 245 26067 430 26079
rect 245 26041 322 26067
rect 245 26007 320 26041
rect 356 26033 430 26067
rect 354 26007 430 26033
rect 245 25999 430 26007
rect 245 25969 322 25999
rect 245 25935 320 25969
rect 356 25965 430 25999
rect 354 25935 430 25965
rect 245 25931 430 25935
rect 245 25897 322 25931
rect 356 25897 430 25931
rect 245 25863 320 25897
rect 354 25863 430 25897
rect 245 25829 322 25863
rect 356 25829 430 25863
rect 245 25825 430 25829
rect 245 25791 320 25825
rect 354 25795 430 25825
rect 245 25761 322 25791
rect 356 25761 430 25795
rect 245 25753 430 25761
rect 245 25719 320 25753
rect 354 25727 430 25753
rect 245 25693 322 25719
rect 356 25693 430 25727
rect 245 25681 430 25693
rect 245 25647 320 25681
rect 354 25659 430 25681
rect 245 25625 322 25647
rect 356 25625 430 25659
rect 245 25609 430 25625
rect 245 25575 320 25609
rect 354 25591 430 25609
rect 245 25557 322 25575
rect 356 25557 430 25591
rect 245 25537 430 25557
rect 245 25503 320 25537
rect 354 25523 430 25537
rect 245 25489 322 25503
rect 356 25489 430 25523
rect 245 25465 430 25489
rect 245 25431 320 25465
rect 354 25455 430 25465
rect 245 25421 322 25431
rect 356 25421 430 25455
rect 245 25393 430 25421
rect 245 25359 320 25393
rect 354 25387 430 25393
rect 245 25353 322 25359
rect 356 25353 430 25387
rect 245 25321 430 25353
rect 245 25287 320 25321
rect 354 25319 430 25321
rect 245 25285 322 25287
rect 356 25285 430 25319
rect 245 25251 430 25285
rect 245 25249 322 25251
rect 245 25215 320 25249
rect 356 25217 430 25251
rect 354 25215 430 25217
rect 245 25183 430 25215
rect 245 25177 322 25183
rect 245 25143 320 25177
rect 356 25149 430 25183
rect 354 25143 430 25149
rect 245 25115 430 25143
rect 245 25105 322 25115
rect 245 25071 320 25105
rect 356 25081 430 25115
rect 354 25071 430 25081
rect 245 25047 430 25071
rect 245 25033 322 25047
rect 245 24999 320 25033
rect 356 25013 430 25047
rect 354 24999 430 25013
rect 245 24979 430 24999
rect 245 24961 322 24979
rect 245 24927 320 24961
rect 356 24945 430 24979
rect 354 24927 430 24945
rect 245 24911 430 24927
rect 245 24889 322 24911
rect 245 24855 320 24889
rect 356 24877 430 24911
rect 354 24855 430 24877
rect 245 24843 430 24855
rect 245 24817 322 24843
rect 245 24783 320 24817
rect 356 24809 430 24843
rect 354 24783 430 24809
rect 245 24775 430 24783
rect 245 24745 322 24775
rect 245 24711 320 24745
rect 356 24741 430 24775
rect 354 24711 430 24741
rect 245 24707 430 24711
rect 245 24673 322 24707
rect 356 24673 430 24707
rect 245 24639 320 24673
rect 354 24639 430 24673
rect 245 24605 322 24639
rect 356 24605 430 24639
rect 245 24601 430 24605
rect 245 24567 320 24601
rect 354 24571 430 24601
rect 245 24537 322 24567
rect 356 24537 430 24571
rect 245 24529 430 24537
rect 245 24495 320 24529
rect 354 24503 430 24529
rect 245 24469 322 24495
rect 356 24469 430 24503
rect 245 24457 430 24469
rect 245 24423 320 24457
rect 354 24435 430 24457
rect 245 24401 322 24423
rect 356 24401 430 24435
rect 245 24385 430 24401
rect 245 24351 320 24385
rect 354 24367 430 24385
rect 245 24333 322 24351
rect 356 24333 430 24367
rect 245 24313 430 24333
rect 245 24279 320 24313
rect 354 24299 430 24313
rect 245 24265 322 24279
rect 356 24265 430 24299
rect 245 24241 430 24265
rect 245 24207 320 24241
rect 354 24231 430 24241
rect 245 24197 322 24207
rect 356 24197 430 24231
rect 245 24169 430 24197
rect 245 24135 320 24169
rect 354 24163 430 24169
rect 245 24129 322 24135
rect 356 24129 430 24163
rect 245 24097 430 24129
rect 245 24063 320 24097
rect 354 24095 430 24097
rect 245 24061 322 24063
rect 356 24061 430 24095
rect 245 24027 430 24061
rect 245 24025 322 24027
rect 245 23991 320 24025
rect 356 23993 430 24027
rect 354 23991 430 23993
rect 245 23959 430 23991
rect 245 23953 322 23959
rect 245 23919 320 23953
rect 356 23925 430 23959
rect 354 23919 430 23925
rect 245 23891 430 23919
rect 245 23881 322 23891
rect 245 23847 320 23881
rect 356 23857 430 23891
rect 354 23847 430 23857
rect 245 23823 430 23847
rect 245 23809 322 23823
rect 245 23775 320 23809
rect 356 23789 430 23823
rect 354 23775 430 23789
rect 245 23755 430 23775
rect 245 23737 322 23755
rect 245 23703 320 23737
rect 356 23721 430 23755
rect 354 23703 430 23721
rect 245 23687 430 23703
rect 245 23665 322 23687
rect 245 23631 320 23665
rect 356 23653 430 23687
rect 354 23631 430 23653
rect 245 23619 430 23631
rect 245 23593 322 23619
rect 245 23559 320 23593
rect 356 23585 430 23619
rect 354 23559 430 23585
rect 245 23551 430 23559
rect 245 23521 322 23551
rect 245 23487 320 23521
rect 356 23517 430 23551
rect 354 23487 430 23517
rect 245 23483 430 23487
rect 245 23449 322 23483
rect 356 23449 430 23483
rect 245 23415 320 23449
rect 354 23415 430 23449
rect 245 23381 322 23415
rect 356 23381 430 23415
rect 245 23377 430 23381
rect 245 23343 320 23377
rect 354 23347 430 23377
rect 245 23313 322 23343
rect 356 23313 430 23347
rect 245 23305 430 23313
rect 245 23271 320 23305
rect 354 23279 430 23305
rect 245 23245 322 23271
rect 356 23245 430 23279
rect 245 23233 430 23245
rect 245 23199 320 23233
rect 354 23211 430 23233
rect 245 23177 322 23199
rect 356 23177 430 23211
rect 245 23161 430 23177
rect 245 23127 320 23161
rect 354 23143 430 23161
rect 245 23109 322 23127
rect 356 23109 430 23143
rect 245 23089 430 23109
rect 245 23055 320 23089
rect 354 23075 430 23089
rect 245 23041 322 23055
rect 356 23041 430 23075
rect 245 23017 430 23041
rect 245 22983 320 23017
rect 354 23007 430 23017
rect 245 22973 322 22983
rect 356 22973 430 23007
rect 245 22945 430 22973
rect 245 22911 320 22945
rect 354 22939 430 22945
rect 245 22905 322 22911
rect 356 22905 430 22939
rect 245 22873 430 22905
rect 245 22839 320 22873
rect 354 22871 430 22873
rect 245 22837 322 22839
rect 356 22837 430 22871
rect 245 22803 430 22837
rect 245 22801 322 22803
rect 245 22767 320 22801
rect 356 22769 430 22803
rect 354 22767 430 22769
rect 245 22735 430 22767
rect 245 22729 322 22735
rect 245 22695 320 22729
rect 356 22701 430 22735
rect 354 22695 430 22701
rect 245 22667 430 22695
rect 245 22657 322 22667
rect 245 22623 320 22657
rect 356 22633 430 22667
rect 354 22623 430 22633
rect 245 22599 430 22623
rect 245 22585 322 22599
rect 245 22551 320 22585
rect 356 22565 430 22599
rect 354 22551 430 22565
rect 245 22531 430 22551
rect 245 22513 322 22531
rect 245 22479 320 22513
rect 356 22497 430 22531
rect 354 22479 430 22497
rect 245 22463 430 22479
rect 245 22441 322 22463
rect 245 22407 320 22441
rect 356 22429 430 22463
rect 354 22407 430 22429
rect 245 22395 430 22407
rect 245 22369 322 22395
rect 245 22335 320 22369
rect 356 22361 430 22395
rect 354 22335 430 22361
rect 245 22327 430 22335
rect 245 22297 322 22327
rect 245 22263 320 22297
rect 356 22293 430 22327
rect 354 22263 430 22293
rect 245 22259 430 22263
rect 245 22225 322 22259
rect 356 22225 430 22259
rect 245 22191 320 22225
rect 354 22191 430 22225
rect 245 22157 322 22191
rect 356 22157 430 22191
rect 245 22153 430 22157
rect 245 22119 320 22153
rect 354 22123 430 22153
rect 245 22089 322 22119
rect 356 22089 430 22123
rect 245 22081 430 22089
rect 245 22047 320 22081
rect 354 22055 430 22081
rect 245 22021 322 22047
rect 356 22021 430 22055
rect 245 22009 430 22021
rect 245 21975 320 22009
rect 354 21987 430 22009
rect 245 21953 322 21975
rect 356 21953 430 21987
rect 245 21937 430 21953
rect 245 21903 320 21937
rect 354 21919 430 21937
rect 245 21885 322 21903
rect 356 21885 430 21919
rect 245 21865 430 21885
rect 245 21831 320 21865
rect 354 21851 430 21865
rect 245 21817 322 21831
rect 356 21817 430 21851
rect 245 21793 430 21817
rect 245 21759 320 21793
rect 354 21783 430 21793
rect 245 21749 322 21759
rect 356 21749 430 21783
rect 245 21721 430 21749
rect 245 21687 320 21721
rect 354 21715 430 21721
rect 245 21681 322 21687
rect 356 21681 430 21715
rect 245 21649 430 21681
rect 245 21615 320 21649
rect 354 21647 430 21649
rect 245 21613 322 21615
rect 356 21613 430 21647
rect 245 21579 430 21613
rect 245 21577 322 21579
rect 245 21543 320 21577
rect 356 21545 430 21579
rect 354 21543 430 21545
rect 245 21511 430 21543
rect 245 21505 322 21511
rect 245 21471 320 21505
rect 356 21477 430 21511
rect 354 21471 430 21477
rect 245 21443 430 21471
rect 245 21433 322 21443
rect 245 21399 320 21433
rect 356 21409 430 21443
rect 354 21399 430 21409
rect 245 21375 430 21399
rect 245 21361 322 21375
rect 245 21327 320 21361
rect 356 21341 430 21375
rect 354 21327 430 21341
rect 245 21307 430 21327
rect 245 21289 322 21307
rect 245 21255 320 21289
rect 356 21273 430 21307
rect 354 21255 430 21273
rect 245 21239 430 21255
rect 245 21217 322 21239
rect 245 21183 320 21217
rect 356 21205 430 21239
rect 354 21183 430 21205
rect 245 21171 430 21183
rect 245 21145 322 21171
rect 245 21111 320 21145
rect 356 21137 430 21171
rect 354 21111 430 21137
rect 245 21103 430 21111
rect 245 21073 322 21103
rect 245 21039 320 21073
rect 356 21069 430 21103
rect 354 21039 430 21069
rect 245 21035 430 21039
rect 245 21001 322 21035
rect 356 21001 430 21035
rect 245 20967 320 21001
rect 354 20967 430 21001
rect 245 20933 322 20967
rect 356 20933 430 20967
rect 245 20929 430 20933
rect 245 20895 320 20929
rect 354 20899 430 20929
rect 245 20865 322 20895
rect 356 20865 430 20899
rect 245 20857 430 20865
rect 245 20823 320 20857
rect 354 20831 430 20857
rect 245 20797 322 20823
rect 356 20797 430 20831
rect 245 20785 430 20797
rect 245 20751 320 20785
rect 354 20763 430 20785
rect 245 20729 322 20751
rect 356 20729 430 20763
rect 245 20713 430 20729
rect 245 20679 320 20713
rect 354 20695 430 20713
rect 245 20661 322 20679
rect 356 20661 430 20695
rect 245 20641 430 20661
rect 245 20607 320 20641
rect 354 20627 430 20641
rect 245 20593 322 20607
rect 356 20593 430 20627
rect 245 20569 430 20593
rect 245 20535 320 20569
rect 354 20559 430 20569
rect 245 20525 322 20535
rect 356 20525 430 20559
rect 245 20497 430 20525
rect 245 20463 320 20497
rect 354 20491 430 20497
rect 245 20457 322 20463
rect 356 20457 430 20491
rect 245 20425 430 20457
rect 245 20391 320 20425
rect 354 20423 430 20425
rect 245 20389 322 20391
rect 356 20389 430 20423
rect 245 20355 430 20389
rect 245 20353 322 20355
rect 245 20319 320 20353
rect 356 20321 430 20355
rect 354 20319 430 20321
rect 245 20287 430 20319
rect 245 20281 322 20287
rect 245 20247 320 20281
rect 356 20253 430 20287
rect 354 20247 430 20253
rect 245 20219 430 20247
rect 245 20209 322 20219
rect 245 20175 320 20209
rect 356 20185 430 20219
rect 354 20175 430 20185
rect 245 20151 430 20175
rect 245 20137 322 20151
rect 245 20103 320 20137
rect 356 20117 430 20151
rect 354 20103 430 20117
rect 245 20083 430 20103
rect 245 20065 322 20083
rect 245 20031 320 20065
rect 356 20049 430 20083
rect 354 20031 430 20049
rect 245 20015 430 20031
rect 245 19993 322 20015
rect 245 19959 320 19993
rect 356 19981 430 20015
rect 354 19959 430 19981
rect 245 19947 430 19959
rect 245 19921 322 19947
rect 245 19887 320 19921
rect 356 19913 430 19947
rect 354 19887 430 19913
rect 245 19879 430 19887
rect 245 19849 322 19879
rect 245 19815 320 19849
rect 356 19845 430 19879
rect 354 19815 430 19845
rect 245 19811 430 19815
rect 245 19777 322 19811
rect 356 19777 430 19811
rect 245 19743 320 19777
rect 354 19743 430 19777
rect 245 19709 322 19743
rect 356 19709 430 19743
rect 245 19705 430 19709
rect 245 19671 320 19705
rect 354 19675 430 19705
rect 245 19641 322 19671
rect 356 19641 430 19675
rect 245 19633 430 19641
rect 245 19599 320 19633
rect 354 19607 430 19633
rect 245 19573 322 19599
rect 356 19573 430 19607
rect 245 19561 430 19573
rect 245 19527 320 19561
rect 354 19539 430 19561
rect 245 19505 322 19527
rect 356 19505 430 19539
rect 245 19489 430 19505
rect 245 19455 320 19489
rect 354 19471 430 19489
rect 245 19437 322 19455
rect 356 19437 430 19471
rect 245 19417 430 19437
rect 245 19383 320 19417
rect 354 19403 430 19417
rect 245 19369 322 19383
rect 356 19369 430 19403
rect 245 19345 430 19369
rect 245 19311 320 19345
rect 354 19335 430 19345
rect 245 19301 322 19311
rect 356 19301 430 19335
rect 245 19273 430 19301
rect 245 19239 320 19273
rect 354 19267 430 19273
rect 245 19233 322 19239
rect 356 19233 430 19267
rect 245 19201 430 19233
rect 245 19167 320 19201
rect 354 19199 430 19201
rect 245 19165 322 19167
rect 356 19165 430 19199
rect 245 19131 430 19165
rect 245 19129 322 19131
rect 245 19095 320 19129
rect 356 19097 430 19131
rect 354 19095 430 19097
rect 245 19063 430 19095
rect 245 19057 322 19063
rect 245 19023 320 19057
rect 356 19029 430 19063
rect 354 19023 430 19029
rect 245 18995 430 19023
rect 245 18985 322 18995
rect 245 18951 320 18985
rect 356 18961 430 18995
rect 354 18951 430 18961
rect 245 18927 430 18951
rect 245 18913 322 18927
rect 245 18879 320 18913
rect 356 18893 430 18927
rect 354 18879 430 18893
rect 245 18859 430 18879
rect 245 18841 322 18859
rect 245 18807 320 18841
rect 356 18825 430 18859
rect 354 18807 430 18825
rect 245 18791 430 18807
rect 245 18769 322 18791
rect 245 18735 320 18769
rect 356 18757 430 18791
rect 354 18735 430 18757
rect 245 18723 430 18735
rect 245 18697 322 18723
rect 245 18663 320 18697
rect 356 18689 430 18723
rect 354 18663 430 18689
rect 245 18655 430 18663
rect 245 18625 322 18655
rect 245 18591 320 18625
rect 356 18621 430 18655
rect 354 18591 430 18621
rect 245 18587 430 18591
rect 245 18553 322 18587
rect 356 18553 430 18587
rect 245 18519 320 18553
rect 354 18519 430 18553
rect 245 18485 322 18519
rect 356 18485 430 18519
rect 245 18481 430 18485
rect 245 18447 320 18481
rect 354 18451 430 18481
rect 245 18417 322 18447
rect 356 18417 430 18451
rect 245 18409 430 18417
rect 245 18375 320 18409
rect 354 18383 430 18409
rect 245 18349 322 18375
rect 356 18349 430 18383
rect 245 18337 430 18349
rect 245 18303 320 18337
rect 354 18315 430 18337
rect 245 18281 322 18303
rect 356 18281 430 18315
rect 245 18265 430 18281
rect 245 18231 320 18265
rect 354 18247 430 18265
rect 245 18213 322 18231
rect 356 18213 430 18247
rect 245 18193 430 18213
rect 245 18159 320 18193
rect 354 18179 430 18193
rect 245 18145 322 18159
rect 356 18145 430 18179
rect 245 18121 430 18145
rect 245 18087 320 18121
rect 354 18111 430 18121
rect 245 18077 322 18087
rect 356 18077 430 18111
rect 245 18049 430 18077
rect 245 18015 320 18049
rect 354 18043 430 18049
rect 245 18009 322 18015
rect 356 18009 430 18043
rect 245 17977 430 18009
rect 245 17943 320 17977
rect 354 17975 430 17977
rect 245 17941 322 17943
rect 356 17941 430 17975
rect 245 17907 430 17941
rect 245 17905 322 17907
rect 245 17871 320 17905
rect 356 17873 430 17907
rect 354 17871 430 17873
rect 245 17839 430 17871
rect 245 17833 322 17839
rect 245 17799 320 17833
rect 356 17805 430 17839
rect 354 17799 430 17805
rect 245 17771 430 17799
rect 245 17761 322 17771
rect 245 17727 320 17761
rect 356 17737 430 17771
rect 354 17727 430 17737
rect 245 17703 430 17727
rect 245 17689 322 17703
rect 245 17655 320 17689
rect 356 17669 430 17703
rect 354 17655 430 17669
rect 245 17635 430 17655
rect 245 17617 322 17635
rect 245 17583 320 17617
rect 356 17601 430 17635
rect 354 17583 430 17601
rect 245 17567 430 17583
rect 245 17545 322 17567
rect 245 17511 320 17545
rect 356 17533 430 17567
rect 354 17511 430 17533
rect 245 17499 430 17511
rect 245 17473 322 17499
rect 245 17439 320 17473
rect 356 17465 430 17499
rect 354 17439 430 17465
rect 245 17431 430 17439
rect 245 17401 322 17431
rect 245 17367 320 17401
rect 356 17397 430 17431
rect 354 17367 430 17397
rect 245 17363 430 17367
rect 245 17329 322 17363
rect 356 17329 430 17363
rect 245 17295 320 17329
rect 354 17295 430 17329
rect 245 17261 322 17295
rect 356 17261 430 17295
rect 245 17257 430 17261
rect 245 17223 320 17257
rect 354 17227 430 17257
rect 245 17193 322 17223
rect 356 17193 430 17227
rect 245 17185 430 17193
rect 245 17151 320 17185
rect 354 17159 430 17185
rect 245 17125 322 17151
rect 356 17125 430 17159
rect 245 17113 430 17125
rect 245 17079 320 17113
rect 354 17091 430 17113
rect 245 17057 322 17079
rect 356 17057 430 17091
rect 245 17041 430 17057
rect 245 17007 320 17041
rect 354 17023 430 17041
rect 245 16989 322 17007
rect 356 16989 430 17023
rect 245 16969 430 16989
rect 245 16935 320 16969
rect 354 16955 430 16969
rect 245 16921 322 16935
rect 356 16921 430 16955
rect 245 16897 430 16921
rect 245 16863 320 16897
rect 354 16887 430 16897
rect 245 16853 322 16863
rect 356 16853 430 16887
rect 245 16825 430 16853
rect 245 16791 320 16825
rect 354 16819 430 16825
rect 245 16785 322 16791
rect 356 16785 430 16819
rect 245 16753 430 16785
rect 245 16719 320 16753
rect 354 16751 430 16753
rect 245 16717 322 16719
rect 356 16717 430 16751
rect 245 16683 430 16717
rect 245 16681 322 16683
rect 245 16647 320 16681
rect 356 16649 430 16683
rect 354 16647 430 16649
rect 245 16615 430 16647
rect 245 16609 322 16615
rect 245 16575 320 16609
rect 356 16581 430 16615
rect 354 16575 430 16581
rect 245 16547 430 16575
rect 245 16537 322 16547
rect 245 16503 320 16537
rect 356 16513 430 16547
rect 354 16503 430 16513
rect 245 16479 430 16503
rect 245 16465 322 16479
rect 245 16431 320 16465
rect 356 16445 430 16479
rect 354 16431 430 16445
rect 245 16411 430 16431
rect 245 16393 322 16411
rect 245 16359 320 16393
rect 356 16377 430 16411
rect 354 16359 430 16377
rect 245 16343 430 16359
rect 245 16321 322 16343
rect 245 16287 320 16321
rect 356 16309 430 16343
rect 354 16287 430 16309
rect 245 16275 430 16287
rect 245 16249 322 16275
rect 245 16215 320 16249
rect 356 16241 430 16275
rect 354 16215 430 16241
rect 245 16207 430 16215
rect 245 16177 322 16207
rect 245 16143 320 16177
rect 356 16173 430 16207
rect 354 16143 430 16173
rect 245 16139 430 16143
rect 245 16105 322 16139
rect 356 16105 430 16139
rect 245 16071 320 16105
rect 354 16071 430 16105
rect 245 16037 322 16071
rect 356 16037 430 16071
rect 245 16033 430 16037
rect 245 15999 320 16033
rect 354 16003 430 16033
rect 245 15969 322 15999
rect 356 15969 430 16003
rect 245 15961 430 15969
rect 245 15927 320 15961
rect 354 15935 430 15961
rect 245 15901 322 15927
rect 356 15901 430 15935
rect 245 15889 430 15901
rect 245 15855 320 15889
rect 354 15867 430 15889
rect 245 15833 322 15855
rect 356 15833 430 15867
rect 245 15817 430 15833
rect 245 15783 320 15817
rect 354 15799 430 15817
rect 245 15765 322 15783
rect 356 15765 430 15799
rect 245 15745 430 15765
rect 245 15711 320 15745
rect 354 15731 430 15745
rect 245 15697 322 15711
rect 356 15697 430 15731
rect 245 15673 430 15697
rect 245 15639 320 15673
rect 354 15663 430 15673
rect 245 15629 322 15639
rect 356 15629 430 15663
rect 245 15601 430 15629
rect 245 15567 320 15601
rect 354 15595 430 15601
rect 245 15561 322 15567
rect 356 15561 430 15595
rect 245 15529 430 15561
rect 245 15495 320 15529
rect 354 15527 430 15529
rect 245 15493 322 15495
rect 356 15493 430 15527
rect 245 15459 430 15493
rect 245 15457 322 15459
rect 245 15423 320 15457
rect 356 15425 430 15459
rect 354 15423 430 15425
rect 245 15391 430 15423
rect 245 15385 322 15391
rect 245 15351 320 15385
rect 356 15357 430 15391
rect 354 15351 430 15357
rect 245 15323 430 15351
rect 245 15313 322 15323
rect 245 15279 320 15313
rect 356 15289 430 15323
rect 354 15279 430 15289
rect 245 15255 430 15279
rect 245 15241 322 15255
rect 245 15207 320 15241
rect 356 15221 430 15255
rect 354 15207 430 15221
rect 245 15187 430 15207
rect 245 15169 322 15187
rect 245 15135 320 15169
rect 356 15153 430 15187
rect 354 15135 430 15153
rect 245 15119 430 15135
rect 245 15097 322 15119
rect 245 15063 320 15097
rect 356 15085 430 15119
rect 354 15063 430 15085
rect 245 15051 430 15063
rect 245 15025 322 15051
rect 245 14991 320 15025
rect 356 15017 430 15051
rect 354 14991 430 15017
rect 245 14983 430 14991
rect 245 14953 322 14983
rect 245 14919 320 14953
rect 356 14949 430 14983
rect 354 14919 430 14949
rect 245 14915 430 14919
rect 245 14881 322 14915
rect 356 14881 430 14915
rect 245 14847 320 14881
rect 354 14847 430 14881
rect 245 14813 322 14847
rect 356 14813 430 14847
rect 245 14809 430 14813
rect 245 14775 320 14809
rect 354 14779 430 14809
rect 245 14745 322 14775
rect 356 14745 430 14779
rect 245 14737 430 14745
rect 245 14703 320 14737
rect 354 14711 430 14737
rect 245 14677 322 14703
rect 356 14677 430 14711
rect 245 14665 430 14677
rect 245 14631 320 14665
rect 354 14643 430 14665
rect 245 14609 322 14631
rect 356 14609 430 14643
rect 245 14593 430 14609
rect 245 14559 320 14593
rect 354 14575 430 14593
rect 245 14541 322 14559
rect 356 14541 430 14575
rect 245 14521 430 14541
rect 245 14487 320 14521
rect 354 14507 430 14521
rect 245 14473 322 14487
rect 356 14473 430 14507
rect 245 14449 430 14473
rect 245 14415 320 14449
rect 354 14439 430 14449
rect 245 14405 322 14415
rect 356 14405 430 14439
rect 245 14377 430 14405
rect 245 14343 320 14377
rect 354 14371 430 14377
rect 245 14337 322 14343
rect 356 14337 430 14371
rect 245 14305 430 14337
rect 245 14271 320 14305
rect 354 14303 430 14305
rect 245 14269 322 14271
rect 356 14269 430 14303
rect 245 14235 430 14269
rect 245 14233 322 14235
rect 245 14199 320 14233
rect 356 14201 430 14235
rect 354 14199 430 14201
rect 245 14167 430 14199
rect 245 14161 322 14167
rect 245 14127 320 14161
rect 356 14133 430 14167
rect 354 14127 430 14133
rect 245 14099 430 14127
rect 245 14089 322 14099
rect 245 14055 320 14089
rect 356 14065 430 14099
rect 354 14055 430 14065
rect 245 14031 430 14055
rect 245 14017 322 14031
rect 245 13983 320 14017
rect 356 13997 430 14031
rect 354 13983 430 13997
rect 245 13963 430 13983
rect 245 13945 322 13963
rect 245 13911 320 13945
rect 356 13929 430 13963
rect 354 13911 430 13929
rect 245 13895 430 13911
rect 245 13873 322 13895
rect 245 13839 320 13873
rect 356 13861 430 13895
rect 354 13839 430 13861
rect 245 13827 430 13839
rect 245 13801 322 13827
rect 245 13767 320 13801
rect 356 13793 430 13827
rect 354 13767 430 13793
rect 245 13759 430 13767
rect 245 13729 322 13759
rect 245 13695 320 13729
rect 356 13725 430 13759
rect 354 13695 430 13725
rect 245 13691 430 13695
rect 245 13657 322 13691
rect 356 13657 430 13691
rect 245 13623 320 13657
rect 354 13623 430 13657
rect 245 13589 322 13623
rect 356 13589 430 13623
rect 245 13585 430 13589
rect 245 13551 320 13585
rect 354 13555 430 13585
rect 245 13521 322 13551
rect 356 13521 430 13555
rect 245 13513 430 13521
rect 245 13479 320 13513
rect 354 13487 430 13513
rect 245 13453 322 13479
rect 356 13453 430 13487
rect 245 13441 430 13453
rect 245 13407 320 13441
rect 354 13419 430 13441
rect 245 13385 322 13407
rect 356 13385 430 13419
rect 245 13369 430 13385
rect 245 13335 320 13369
rect 354 13351 430 13369
rect 245 13317 322 13335
rect 356 13317 430 13351
rect 245 13297 430 13317
rect 245 13263 320 13297
rect 354 13283 430 13297
rect 245 13249 322 13263
rect 356 13249 430 13283
rect 245 13225 430 13249
rect 245 13191 320 13225
rect 354 13215 430 13225
rect 245 13181 322 13191
rect 356 13181 430 13215
rect 245 13153 430 13181
rect 245 13119 320 13153
rect 354 13147 430 13153
rect 245 13113 322 13119
rect 356 13113 430 13147
rect 245 13081 430 13113
rect 245 13047 320 13081
rect 354 13079 430 13081
rect 245 13045 322 13047
rect 356 13045 430 13079
rect 245 13011 430 13045
rect 245 13009 322 13011
rect 245 12975 320 13009
rect 356 12977 430 13011
rect 354 12975 430 12977
rect 245 12943 430 12975
rect 245 12937 322 12943
rect 245 12903 320 12937
rect 356 12909 430 12943
rect 354 12903 430 12909
rect 245 12875 430 12903
rect 245 12865 322 12875
rect 245 12831 320 12865
rect 356 12841 430 12875
rect 354 12831 430 12841
rect 245 12807 430 12831
rect 245 12793 322 12807
rect 245 12759 320 12793
rect 356 12773 430 12807
rect 354 12759 430 12773
rect 245 12739 430 12759
rect 245 12721 322 12739
rect 245 12687 320 12721
rect 356 12705 430 12739
rect 354 12687 430 12705
rect 245 12671 430 12687
rect 245 12649 322 12671
rect 245 12615 320 12649
rect 356 12637 430 12671
rect 354 12615 430 12637
rect 245 12603 430 12615
rect 245 12577 322 12603
rect 245 12543 320 12577
rect 356 12569 430 12603
rect 354 12543 430 12569
rect 245 12535 430 12543
rect 245 12505 322 12535
rect 245 12471 320 12505
rect 356 12501 430 12535
rect 354 12471 430 12501
rect 245 12467 430 12471
rect 245 12433 322 12467
rect 356 12433 430 12467
rect 245 12399 320 12433
rect 354 12399 430 12433
rect 245 12365 322 12399
rect 356 12365 430 12399
rect 245 12361 430 12365
rect 245 12327 320 12361
rect 354 12331 430 12361
rect 245 12297 322 12327
rect 356 12297 430 12331
rect 245 12289 430 12297
rect 245 12255 320 12289
rect 354 12263 430 12289
rect 245 12229 322 12255
rect 356 12229 430 12263
rect 245 12217 430 12229
rect 245 12183 320 12217
rect 354 12195 430 12217
rect 245 12161 322 12183
rect 356 12161 430 12195
rect 245 12145 430 12161
rect 245 12111 320 12145
rect 354 12127 430 12145
rect 245 12093 322 12111
rect 356 12093 430 12127
rect 245 12073 430 12093
rect 245 12039 320 12073
rect 354 12059 430 12073
rect 245 12025 322 12039
rect 356 12025 430 12059
rect 245 12001 430 12025
rect 245 11967 320 12001
rect 354 11991 430 12001
rect 245 11957 322 11967
rect 356 11957 430 11991
rect 245 11929 430 11957
rect 245 11895 320 11929
rect 354 11923 430 11929
rect 245 11889 322 11895
rect 356 11889 430 11923
rect 245 11857 430 11889
rect 245 11823 320 11857
rect 354 11855 430 11857
rect 245 11821 322 11823
rect 356 11821 430 11855
rect 245 11787 430 11821
rect 245 11785 322 11787
rect 245 11751 320 11785
rect 356 11753 430 11787
rect 354 11751 430 11753
rect 245 11719 430 11751
rect 245 11713 322 11719
rect 245 11679 320 11713
rect 356 11685 430 11719
rect 354 11679 430 11685
rect 245 11651 430 11679
rect 245 11641 322 11651
rect 245 11607 320 11641
rect 356 11617 430 11651
rect 354 11607 430 11617
rect 245 11583 430 11607
rect 245 11569 322 11583
rect 245 11535 320 11569
rect 356 11549 430 11583
rect 354 11535 430 11549
rect 245 11515 430 11535
rect 245 11497 322 11515
rect 245 11463 320 11497
rect 356 11481 430 11515
rect 354 11463 430 11481
rect 245 11447 430 11463
rect 245 11425 322 11447
rect 245 11391 320 11425
rect 356 11413 430 11447
rect 354 11391 430 11413
rect 245 11379 430 11391
rect 245 11353 322 11379
rect 245 11319 320 11353
rect 356 11345 430 11379
rect 354 11319 430 11345
rect 245 11311 430 11319
rect 245 11281 322 11311
rect 245 11247 320 11281
rect 356 11277 430 11311
rect 354 11247 430 11277
rect 245 11243 430 11247
rect 245 11209 322 11243
rect 356 11209 430 11243
rect 245 11175 320 11209
rect 354 11175 430 11209
rect 245 11141 322 11175
rect 356 11141 430 11175
rect 245 11137 430 11141
rect 245 11103 320 11137
rect 354 11107 430 11137
rect 245 11073 322 11103
rect 356 11073 430 11107
rect 245 11065 430 11073
rect 245 11031 320 11065
rect 354 11039 430 11065
rect 245 11005 322 11031
rect 356 11005 430 11039
rect 245 10993 430 11005
rect 245 10959 320 10993
rect 354 10971 430 10993
rect 245 10937 322 10959
rect 356 10937 430 10971
rect 245 10921 430 10937
rect 245 10887 320 10921
rect 354 10903 430 10921
rect 245 10869 322 10887
rect 356 10869 430 10903
rect 245 10849 430 10869
rect 245 10815 320 10849
rect 354 10835 430 10849
rect 245 10801 322 10815
rect 356 10801 430 10835
rect 245 10777 430 10801
rect 245 10743 320 10777
rect 354 10767 430 10777
rect 245 10733 322 10743
rect 356 10733 430 10767
rect 245 10705 430 10733
rect 245 10671 320 10705
rect 354 10699 430 10705
rect 245 10665 322 10671
rect 356 10665 430 10699
rect 245 10633 430 10665
rect 245 10599 320 10633
rect 354 10631 430 10633
rect 245 10597 322 10599
rect 356 10597 430 10631
rect 245 10563 430 10597
rect 245 10561 322 10563
rect 245 10527 320 10561
rect 356 10529 430 10563
rect 354 10527 430 10529
rect 245 10495 430 10527
rect 245 10489 322 10495
rect 245 10455 320 10489
rect 356 10461 430 10495
rect 354 10455 430 10461
rect 245 10427 430 10455
rect 245 10417 322 10427
rect 245 10383 320 10417
rect 356 10393 430 10427
rect 354 10383 430 10393
rect 245 10359 430 10383
rect 245 10345 322 10359
rect 245 10311 320 10345
rect 356 10325 430 10359
rect 354 10311 430 10325
rect 245 10291 430 10311
rect 245 10273 322 10291
rect 245 10239 320 10273
rect 356 10257 430 10291
rect 354 10239 430 10257
rect 245 10223 430 10239
rect 245 10201 322 10223
rect 245 10167 320 10201
rect 356 10189 430 10223
rect 354 10167 430 10189
rect 245 10155 430 10167
rect 245 10129 322 10155
rect 245 10095 320 10129
rect 356 10121 430 10155
rect 354 10095 430 10121
rect 245 10087 430 10095
rect 245 10057 322 10087
rect 245 10023 320 10057
rect 356 10053 430 10087
rect 354 10023 430 10053
rect 245 10019 430 10023
rect 245 9985 322 10019
rect 356 9985 430 10019
rect 245 9951 320 9985
rect 354 9951 430 9985
rect 245 9917 322 9951
rect 356 9917 430 9951
rect 245 9913 430 9917
rect 245 9879 320 9913
rect 354 9883 430 9913
rect 245 9849 322 9879
rect 356 9849 430 9883
rect 245 9841 430 9849
rect 245 9807 320 9841
rect 354 9815 430 9841
rect 245 9781 322 9807
rect 356 9781 430 9815
rect 245 9769 430 9781
rect 245 9735 320 9769
rect 354 9747 430 9769
rect 245 9713 322 9735
rect 356 9713 430 9747
rect 245 9697 430 9713
rect 617 36177 14361 36207
rect 617 36143 773 36177
rect 807 36143 841 36177
rect 875 36143 909 36177
rect 943 36143 977 36177
rect 1011 36143 1045 36177
rect 1079 36143 1113 36177
rect 1147 36143 1181 36177
rect 1215 36143 1249 36177
rect 1283 36143 1317 36177
rect 1351 36143 1385 36177
rect 1419 36143 1453 36177
rect 1487 36143 1521 36177
rect 1555 36143 1589 36177
rect 1623 36143 1657 36177
rect 1691 36143 1725 36177
rect 1759 36143 1793 36177
rect 1827 36143 1861 36177
rect 1895 36143 1929 36177
rect 1963 36143 1997 36177
rect 2031 36143 2065 36177
rect 2099 36143 2133 36177
rect 2167 36143 2201 36177
rect 2235 36143 2269 36177
rect 2303 36143 2337 36177
rect 2371 36143 2405 36177
rect 2439 36143 2473 36177
rect 2507 36143 2541 36177
rect 2575 36143 2609 36177
rect 2643 36143 2677 36177
rect 2711 36143 2745 36177
rect 2779 36143 2813 36177
rect 2847 36143 2881 36177
rect 2915 36143 2949 36177
rect 2983 36143 3017 36177
rect 3051 36143 3085 36177
rect 3119 36143 3153 36177
rect 3187 36143 3221 36177
rect 3255 36143 3289 36177
rect 3323 36143 3357 36177
rect 3391 36143 3425 36177
rect 3459 36143 3493 36177
rect 3527 36143 3561 36177
rect 3595 36143 3629 36177
rect 3663 36143 3697 36177
rect 3731 36143 3765 36177
rect 3799 36143 3833 36177
rect 3867 36143 3901 36177
rect 3935 36143 3969 36177
rect 4003 36143 4037 36177
rect 4071 36143 4105 36177
rect 4139 36143 4173 36177
rect 4207 36143 4241 36177
rect 4275 36143 4309 36177
rect 4343 36143 4377 36177
rect 4411 36143 4445 36177
rect 4479 36143 4513 36177
rect 4547 36143 4581 36177
rect 4615 36143 4649 36177
rect 4683 36143 4717 36177
rect 4751 36143 4785 36177
rect 4819 36143 4853 36177
rect 4887 36143 4921 36177
rect 4955 36143 4989 36177
rect 5023 36143 5057 36177
rect 5091 36143 5125 36177
rect 5159 36143 5193 36177
rect 5227 36143 5261 36177
rect 5295 36143 5329 36177
rect 5363 36143 5397 36177
rect 5431 36143 5465 36177
rect 5499 36143 5533 36177
rect 5567 36143 5601 36177
rect 5635 36143 5669 36177
rect 5703 36143 5737 36177
rect 5771 36143 5805 36177
rect 5839 36143 5873 36177
rect 5907 36143 5941 36177
rect 5975 36143 6009 36177
rect 6043 36143 6077 36177
rect 6111 36143 6145 36177
rect 6179 36143 6213 36177
rect 6247 36143 6281 36177
rect 6315 36143 6349 36177
rect 6383 36143 6417 36177
rect 6451 36143 6485 36177
rect 6519 36143 6553 36177
rect 6587 36143 6621 36177
rect 6655 36143 6689 36177
rect 6723 36143 6757 36177
rect 6791 36143 6825 36177
rect 6859 36143 6893 36177
rect 6927 36143 6961 36177
rect 6995 36143 7029 36177
rect 7063 36143 7097 36177
rect 7131 36143 7165 36177
rect 7199 36143 7233 36177
rect 7267 36143 7301 36177
rect 7335 36143 7369 36177
rect 7403 36143 7437 36177
rect 7471 36143 7505 36177
rect 7539 36143 7573 36177
rect 7607 36143 7641 36177
rect 7675 36143 7709 36177
rect 7743 36143 7777 36177
rect 7811 36143 7845 36177
rect 7879 36143 7913 36177
rect 7947 36143 7981 36177
rect 8015 36143 8049 36177
rect 8083 36143 8117 36177
rect 8151 36143 8185 36177
rect 8219 36143 8253 36177
rect 8287 36143 8321 36177
rect 8355 36143 8389 36177
rect 8423 36143 8457 36177
rect 8491 36143 8525 36177
rect 8559 36143 8593 36177
rect 8627 36143 8661 36177
rect 8695 36143 8729 36177
rect 8763 36143 8797 36177
rect 8831 36143 8865 36177
rect 8899 36143 8933 36177
rect 8967 36143 9001 36177
rect 9035 36143 9069 36177
rect 9103 36143 9137 36177
rect 9171 36143 9205 36177
rect 9239 36143 9273 36177
rect 9307 36143 9341 36177
rect 9375 36143 9409 36177
rect 9443 36143 9477 36177
rect 9511 36143 9545 36177
rect 9579 36143 9613 36177
rect 9647 36143 9681 36177
rect 9715 36143 9749 36177
rect 9783 36143 9817 36177
rect 9851 36143 9885 36177
rect 9919 36143 9953 36177
rect 9987 36143 10021 36177
rect 10055 36143 10089 36177
rect 10123 36143 10157 36177
rect 10191 36143 10225 36177
rect 10259 36143 10293 36177
rect 10327 36143 10361 36177
rect 10395 36143 10429 36177
rect 10463 36143 10497 36177
rect 10531 36143 10565 36177
rect 10599 36143 10633 36177
rect 10667 36143 10701 36177
rect 10735 36143 10769 36177
rect 10803 36143 10837 36177
rect 10871 36143 10905 36177
rect 10939 36143 10973 36177
rect 11007 36143 11041 36177
rect 11075 36143 11109 36177
rect 11143 36143 11177 36177
rect 11211 36143 11245 36177
rect 11279 36143 11313 36177
rect 11347 36143 11381 36177
rect 11415 36143 11449 36177
rect 11483 36143 11517 36177
rect 11551 36143 11585 36177
rect 11619 36143 11653 36177
rect 11687 36143 11721 36177
rect 11755 36143 11789 36177
rect 11823 36143 11857 36177
rect 11891 36143 11925 36177
rect 11959 36143 11993 36177
rect 12027 36143 12061 36177
rect 12095 36143 12129 36177
rect 12163 36143 12197 36177
rect 12231 36143 12265 36177
rect 12299 36143 12333 36177
rect 12367 36143 12401 36177
rect 12435 36143 12469 36177
rect 12503 36143 12537 36177
rect 12571 36143 12605 36177
rect 12639 36143 12673 36177
rect 12707 36143 12741 36177
rect 12775 36143 12809 36177
rect 12843 36143 12877 36177
rect 12911 36143 12945 36177
rect 12979 36143 13013 36177
rect 13047 36143 13081 36177
rect 13115 36143 13149 36177
rect 13183 36143 13217 36177
rect 13251 36143 13285 36177
rect 13319 36143 13353 36177
rect 13387 36143 13421 36177
rect 13455 36143 13489 36177
rect 13523 36143 13557 36177
rect 13591 36143 13625 36177
rect 13659 36143 13693 36177
rect 13727 36143 13761 36177
rect 13795 36143 13829 36177
rect 13863 36143 13897 36177
rect 13931 36143 13965 36177
rect 13999 36143 14033 36177
rect 14067 36143 14101 36177
rect 14135 36143 14169 36177
rect 14203 36143 14361 36177
rect 617 36032 14361 36143
rect 617 35998 646 36032
rect 680 36003 14297 36032
rect 680 35998 1009 36003
rect 617 35969 1009 35998
rect 1043 35969 1081 36003
rect 1115 35969 1153 36003
rect 1187 35969 1225 36003
rect 1259 35969 1297 36003
rect 1331 35969 1369 36003
rect 1403 35969 1441 36003
rect 1475 35969 1513 36003
rect 1547 35969 1585 36003
rect 1619 35969 1657 36003
rect 1691 35969 1729 36003
rect 1763 35969 1801 36003
rect 1835 35969 1873 36003
rect 1907 35969 1945 36003
rect 1979 35969 2017 36003
rect 2051 35969 2089 36003
rect 2123 35969 2161 36003
rect 2195 35969 2233 36003
rect 2267 35969 2305 36003
rect 2339 35969 2377 36003
rect 2411 35969 2449 36003
rect 2483 35969 2521 36003
rect 2555 35969 2593 36003
rect 2627 35969 2665 36003
rect 2699 35969 2737 36003
rect 2771 35969 2809 36003
rect 2843 35969 2881 36003
rect 2915 35969 2953 36003
rect 2987 35969 3025 36003
rect 3059 35969 3097 36003
rect 3131 35969 3169 36003
rect 3203 35969 3241 36003
rect 3275 35969 3313 36003
rect 3347 35969 3385 36003
rect 3419 35969 3457 36003
rect 3491 35969 3529 36003
rect 3563 35969 3601 36003
rect 3635 35969 3673 36003
rect 3707 35969 3745 36003
rect 3779 35969 3817 36003
rect 3851 35969 3889 36003
rect 3923 35969 3961 36003
rect 3995 35969 4033 36003
rect 4067 35969 4105 36003
rect 4139 35969 4177 36003
rect 4211 35969 4249 36003
rect 4283 35969 4321 36003
rect 4355 35969 4393 36003
rect 4427 35969 4465 36003
rect 4499 35969 4537 36003
rect 4571 35969 4609 36003
rect 4643 35969 4681 36003
rect 4715 35969 4753 36003
rect 4787 35969 4825 36003
rect 4859 35969 4897 36003
rect 4931 35969 4969 36003
rect 5003 35969 5041 36003
rect 5075 35969 5113 36003
rect 5147 35969 5185 36003
rect 5219 35969 5257 36003
rect 5291 35969 5329 36003
rect 5363 35969 5401 36003
rect 5435 35969 5473 36003
rect 5507 35969 5545 36003
rect 5579 35969 5617 36003
rect 5651 35969 5689 36003
rect 5723 35969 5761 36003
rect 5795 35969 5833 36003
rect 5867 35969 5905 36003
rect 5939 35969 5977 36003
rect 6011 35969 6049 36003
rect 6083 35969 6121 36003
rect 6155 35969 6193 36003
rect 6227 35969 6265 36003
rect 6299 35969 6337 36003
rect 6371 35969 6409 36003
rect 6443 35969 6481 36003
rect 6515 35969 6553 36003
rect 6587 35969 6625 36003
rect 6659 35969 6697 36003
rect 6731 35969 6769 36003
rect 6803 35969 6841 36003
rect 6875 35969 6913 36003
rect 6947 35969 6985 36003
rect 7019 35969 7057 36003
rect 7091 35969 7129 36003
rect 7163 35969 7201 36003
rect 7235 35969 7273 36003
rect 7307 35969 7345 36003
rect 7379 35969 7417 36003
rect 7451 35969 7489 36003
rect 7523 35969 7561 36003
rect 7595 35969 7633 36003
rect 7667 35969 7705 36003
rect 7739 35969 7777 36003
rect 7811 35969 7849 36003
rect 7883 35969 7921 36003
rect 7955 35969 7993 36003
rect 8027 35969 8065 36003
rect 8099 35969 8137 36003
rect 8171 35969 8209 36003
rect 8243 35969 8281 36003
rect 8315 35969 8353 36003
rect 8387 35969 8425 36003
rect 8459 35969 8497 36003
rect 8531 35969 8569 36003
rect 8603 35969 8641 36003
rect 8675 35969 8713 36003
rect 8747 35969 8785 36003
rect 8819 35969 8857 36003
rect 8891 35969 8929 36003
rect 8963 35969 9001 36003
rect 9035 35969 9073 36003
rect 9107 35969 9145 36003
rect 9179 35969 9217 36003
rect 9251 35969 9289 36003
rect 9323 35969 9361 36003
rect 9395 35969 9433 36003
rect 9467 35969 9505 36003
rect 9539 35969 9577 36003
rect 9611 35969 9649 36003
rect 9683 35969 9721 36003
rect 9755 35969 9793 36003
rect 9827 35969 9865 36003
rect 9899 35969 9937 36003
rect 9971 35969 10009 36003
rect 10043 35969 10081 36003
rect 10115 35969 10153 36003
rect 10187 35969 10225 36003
rect 10259 35969 10297 36003
rect 10331 35969 10369 36003
rect 10403 35969 10441 36003
rect 10475 35969 10513 36003
rect 10547 35969 10585 36003
rect 10619 35969 10657 36003
rect 10691 35969 10729 36003
rect 10763 35969 10801 36003
rect 10835 35969 10873 36003
rect 10907 35969 10945 36003
rect 10979 35969 11017 36003
rect 11051 35969 11089 36003
rect 11123 35969 11161 36003
rect 11195 35969 11233 36003
rect 11267 35969 11305 36003
rect 11339 35969 11377 36003
rect 11411 35969 11449 36003
rect 11483 35969 11521 36003
rect 11555 35969 11593 36003
rect 11627 35969 11665 36003
rect 11699 35969 11737 36003
rect 11771 35969 11809 36003
rect 11843 35969 11881 36003
rect 11915 35969 11953 36003
rect 11987 35969 12025 36003
rect 12059 35969 12097 36003
rect 12131 35969 12169 36003
rect 12203 35969 12241 36003
rect 12275 35969 12313 36003
rect 12347 35969 12385 36003
rect 12419 35969 12457 36003
rect 12491 35969 12529 36003
rect 12563 35969 12601 36003
rect 12635 35969 12673 36003
rect 12707 35969 12745 36003
rect 12779 35969 12817 36003
rect 12851 35969 12889 36003
rect 12923 35969 12961 36003
rect 12995 35969 13033 36003
rect 13067 35969 13105 36003
rect 13139 35969 13177 36003
rect 13211 35969 13249 36003
rect 13283 35969 13321 36003
rect 13355 35969 13393 36003
rect 13427 35969 13465 36003
rect 13499 35969 13537 36003
rect 13571 35969 13609 36003
rect 13643 35969 13681 36003
rect 13715 35969 13753 36003
rect 13787 35969 13825 36003
rect 13859 35969 13897 36003
rect 13931 35969 13969 36003
rect 14003 35998 14297 36003
rect 14331 35998 14361 36032
rect 14003 35969 14361 35998
rect 617 35964 14361 35969
rect 617 35930 646 35964
rect 680 35930 14297 35964
rect 14331 35930 14361 35964
rect 617 35911 14361 35930
rect 617 35896 814 35911
rect 617 35862 646 35896
rect 680 35877 814 35896
rect 848 35896 14361 35911
rect 848 35877 14297 35896
rect 680 35862 14297 35877
rect 14331 35862 14361 35896
rect 617 35839 14361 35862
rect 617 35828 814 35839
rect 617 35794 646 35828
rect 680 35805 814 35828
rect 848 35832 14361 35839
rect 848 35805 14120 35832
rect 680 35798 14120 35805
rect 14154 35828 14361 35832
rect 14154 35798 14297 35828
rect 680 35794 14297 35798
rect 14331 35794 14361 35828
rect 617 35767 14361 35794
rect 617 35760 814 35767
rect 617 35726 646 35760
rect 680 35733 814 35760
rect 848 35760 14361 35767
rect 848 35733 14120 35760
rect 680 35726 14120 35733
rect 14154 35726 14297 35760
rect 14331 35726 14361 35760
rect 617 35695 14361 35726
rect 617 35692 814 35695
rect 617 35658 646 35692
rect 680 35661 814 35692
rect 848 35692 14361 35695
rect 848 35688 14297 35692
rect 848 35661 14120 35688
rect 680 35658 14120 35661
rect 617 35654 14120 35658
rect 14154 35658 14297 35688
rect 14331 35658 14361 35692
rect 14154 35654 14361 35658
rect 617 35624 14361 35654
rect 617 35590 646 35624
rect 680 35623 14297 35624
rect 680 35590 814 35623
rect 617 35589 814 35590
rect 848 35616 14297 35623
rect 848 35589 14120 35616
rect 617 35582 14120 35589
rect 14154 35590 14297 35616
rect 14331 35590 14361 35624
rect 14154 35582 14361 35590
rect 617 35556 14361 35582
rect 617 35522 646 35556
rect 680 35551 14297 35556
rect 680 35522 814 35551
rect 617 35517 814 35522
rect 848 35544 14297 35551
rect 848 35517 14120 35544
rect 617 35510 14120 35517
rect 14154 35522 14297 35544
rect 14331 35522 14361 35556
rect 14154 35510 14361 35522
rect 617 35488 14361 35510
rect 617 35454 646 35488
rect 680 35479 14297 35488
rect 680 35454 814 35479
rect 617 35445 814 35454
rect 848 35472 14297 35479
rect 848 35445 14120 35472
rect 617 35438 14120 35445
rect 14154 35454 14297 35472
rect 14331 35454 14361 35488
rect 14154 35438 14361 35454
rect 617 35420 14361 35438
rect 617 35386 646 35420
rect 680 35407 14297 35420
rect 680 35386 814 35407
rect 617 35373 814 35386
rect 848 35400 14297 35407
rect 848 35373 14120 35400
rect 617 35366 14120 35373
rect 14154 35386 14297 35400
rect 14331 35386 14361 35420
rect 14154 35366 14361 35386
rect 617 35352 14361 35366
rect 617 35318 646 35352
rect 680 35335 14297 35352
rect 680 35318 814 35335
rect 617 35301 814 35318
rect 848 35328 14297 35335
rect 848 35301 14120 35328
rect 617 35294 14120 35301
rect 14154 35318 14297 35328
rect 14331 35318 14361 35352
rect 14154 35294 14361 35318
rect 617 35284 14361 35294
rect 617 35250 646 35284
rect 680 35263 14297 35284
rect 680 35250 814 35263
rect 617 35229 814 35250
rect 848 35256 14297 35263
rect 848 35229 14120 35256
rect 617 35222 14120 35229
rect 14154 35250 14297 35256
rect 14331 35250 14361 35284
rect 14154 35222 14361 35250
rect 617 35216 14361 35222
rect 617 35182 646 35216
rect 680 35191 14297 35216
rect 680 35182 814 35191
rect 617 35157 814 35182
rect 848 35184 14297 35191
rect 848 35157 14120 35184
rect 617 35150 14120 35157
rect 14154 35182 14297 35184
rect 14331 35182 14361 35216
rect 14154 35150 14361 35182
rect 617 35148 14361 35150
rect 617 35114 646 35148
rect 680 35119 14297 35148
rect 680 35114 814 35119
rect 617 35085 814 35114
rect 848 35114 14297 35119
rect 14331 35114 14361 35148
rect 848 35112 14361 35114
rect 848 35085 14120 35112
rect 617 35080 14120 35085
rect 617 35046 646 35080
rect 680 35078 14120 35080
rect 14154 35080 14361 35112
rect 14154 35078 14297 35080
rect 680 35047 14297 35078
rect 680 35046 814 35047
rect 617 35013 814 35046
rect 848 35046 14297 35047
rect 14331 35046 14361 35080
rect 848 35040 14361 35046
rect 848 35013 14120 35040
rect 617 35012 14120 35013
rect 617 34978 646 35012
rect 680 35006 14120 35012
rect 14154 35012 14361 35040
rect 14154 35006 14297 35012
rect 680 34978 14297 35006
rect 14331 34978 14361 35012
rect 617 34975 14361 34978
rect 617 34944 814 34975
rect 617 34910 646 34944
rect 680 34941 814 34944
rect 848 34968 14361 34975
rect 848 34941 14120 34968
rect 680 34934 14120 34941
rect 14154 34944 14361 34968
rect 14154 34934 14297 34944
rect 680 34910 14297 34934
rect 14331 34910 14361 34944
rect 617 34903 14361 34910
rect 617 34876 814 34903
rect 617 34842 646 34876
rect 680 34869 814 34876
rect 848 34896 14361 34903
rect 848 34869 14120 34896
rect 680 34862 14120 34869
rect 14154 34876 14361 34896
rect 14154 34862 14297 34876
rect 680 34842 14297 34862
rect 14331 34842 14361 34876
rect 617 34831 14361 34842
rect 617 34808 814 34831
rect 617 34774 646 34808
rect 680 34797 814 34808
rect 848 34797 1026 34831
rect 680 34774 1026 34797
rect 617 34759 1026 34774
rect 617 34740 814 34759
rect 617 34706 646 34740
rect 680 34725 814 34740
rect 848 34725 1026 34759
rect 680 34706 1026 34725
rect 617 34687 1026 34706
rect 617 34672 814 34687
rect 617 34638 646 34672
rect 680 34653 814 34672
rect 848 34653 1026 34687
rect 13968 34824 14361 34831
rect 13968 34790 14120 34824
rect 14154 34808 14361 34824
rect 14154 34790 14297 34808
rect 13968 34774 14297 34790
rect 14331 34774 14361 34808
rect 13968 34752 14361 34774
rect 13968 34718 14120 34752
rect 14154 34740 14361 34752
rect 14154 34718 14297 34740
rect 13968 34706 14297 34718
rect 14331 34706 14361 34740
rect 680 34638 1026 34653
rect 617 34615 1026 34638
rect 617 34604 814 34615
rect 617 34570 646 34604
rect 680 34581 814 34604
rect 848 34581 1026 34615
rect 680 34570 1026 34581
rect 617 34543 1026 34570
rect 617 34536 814 34543
rect 617 34502 646 34536
rect 680 34509 814 34536
rect 848 34509 1026 34543
rect 680 34502 1026 34509
rect 617 34471 1026 34502
rect 617 34468 814 34471
rect 617 34434 646 34468
rect 680 34437 814 34468
rect 848 34437 1026 34471
rect 680 34434 1026 34437
rect 617 34400 1026 34434
rect 617 34366 646 34400
rect 680 34399 1026 34400
rect 680 34366 814 34399
rect 617 34365 814 34366
rect 848 34365 1026 34399
rect 617 34332 1026 34365
rect 617 34298 646 34332
rect 680 34327 1026 34332
rect 680 34298 814 34327
rect 617 34293 814 34298
rect 848 34293 1026 34327
rect 617 34264 1026 34293
rect 617 34230 646 34264
rect 680 34255 1026 34264
rect 680 34230 814 34255
rect 617 34221 814 34230
rect 848 34221 1026 34255
rect 617 34196 1026 34221
rect 617 34162 646 34196
rect 680 34183 1026 34196
rect 680 34162 814 34183
rect 617 34149 814 34162
rect 848 34149 1026 34183
rect 617 34128 1026 34149
rect 617 34094 646 34128
rect 680 34111 1026 34128
rect 680 34094 814 34111
rect 617 34077 814 34094
rect 848 34077 1026 34111
rect 617 34060 1026 34077
rect 617 34026 646 34060
rect 680 34039 1026 34060
rect 680 34026 814 34039
rect 617 34005 814 34026
rect 848 34005 1026 34039
rect 617 33992 1026 34005
rect 617 33958 646 33992
rect 680 33967 1026 33992
rect 680 33958 814 33967
rect 617 33933 814 33958
rect 848 33933 1026 33967
rect 617 33924 1026 33933
rect 617 33890 646 33924
rect 680 33895 1026 33924
rect 680 33890 814 33895
rect 617 33861 814 33890
rect 848 33861 1026 33895
rect 617 33856 1026 33861
rect 617 33822 646 33856
rect 680 33823 1026 33856
rect 680 33822 814 33823
rect 617 33789 814 33822
rect 848 33789 1026 33823
rect 617 33788 1026 33789
rect 617 33754 646 33788
rect 680 33754 1026 33788
rect 617 33751 1026 33754
rect 617 33720 814 33751
rect 617 33686 646 33720
rect 680 33717 814 33720
rect 848 33717 1026 33751
rect 680 33686 1026 33717
rect 617 33679 1026 33686
rect 617 33652 814 33679
rect 617 33618 646 33652
rect 680 33645 814 33652
rect 848 33645 1026 33679
rect 680 33618 1026 33645
rect 617 33607 1026 33618
rect 617 33584 814 33607
rect 617 33550 646 33584
rect 680 33573 814 33584
rect 848 33573 1026 33607
rect 680 33550 1026 33573
rect 617 33535 1026 33550
rect 617 33516 814 33535
rect 617 33482 646 33516
rect 680 33501 814 33516
rect 848 33501 1026 33535
rect 680 33482 1026 33501
rect 617 33463 1026 33482
rect 617 33448 814 33463
rect 617 33414 646 33448
rect 680 33429 814 33448
rect 848 33429 1026 33463
rect 680 33414 1026 33429
rect 617 33391 1026 33414
rect 617 33380 814 33391
rect 617 33346 646 33380
rect 680 33357 814 33380
rect 848 33357 1026 33391
rect 680 33346 1026 33357
rect 617 33319 1026 33346
rect 617 33312 814 33319
rect 617 33278 646 33312
rect 680 33285 814 33312
rect 848 33285 1026 33319
rect 680 33278 1026 33285
rect 617 33247 1026 33278
rect 617 33244 814 33247
rect 617 33210 646 33244
rect 680 33213 814 33244
rect 848 33213 1026 33247
rect 680 33210 1026 33213
rect 617 33176 1026 33210
rect 617 33142 646 33176
rect 680 33175 1026 33176
rect 680 33142 814 33175
rect 617 33141 814 33142
rect 848 33141 1026 33175
rect 617 33108 1026 33141
rect 617 33074 646 33108
rect 680 33103 1026 33108
rect 680 33074 814 33103
rect 617 33069 814 33074
rect 848 33069 1026 33103
rect 617 33040 1026 33069
rect 617 33006 646 33040
rect 680 33031 1026 33040
rect 680 33006 814 33031
rect 617 32997 814 33006
rect 848 32997 1026 33031
rect 617 32972 1026 32997
rect 617 32938 646 32972
rect 680 32959 1026 32972
rect 680 32938 814 32959
rect 617 32925 814 32938
rect 848 32925 1026 32959
rect 617 32904 1026 32925
rect 617 32870 646 32904
rect 680 32887 1026 32904
rect 680 32870 814 32887
rect 617 32853 814 32870
rect 848 32853 1026 32887
rect 617 32836 1026 32853
rect 617 32802 646 32836
rect 680 32815 1026 32836
rect 680 32802 814 32815
rect 617 32781 814 32802
rect 848 32781 1026 32815
rect 617 32768 1026 32781
rect 617 32734 646 32768
rect 680 32743 1026 32768
rect 680 32734 814 32743
rect 617 32709 814 32734
rect 848 32709 1026 32743
rect 617 32700 1026 32709
rect 617 32666 646 32700
rect 680 32671 1026 32700
rect 680 32666 814 32671
rect 617 32637 814 32666
rect 848 32637 1026 32671
rect 617 32632 1026 32637
rect 617 32598 646 32632
rect 680 32599 1026 32632
rect 680 32598 814 32599
rect 617 32565 814 32598
rect 848 32565 1026 32599
rect 617 32564 1026 32565
rect 617 32530 646 32564
rect 680 32530 1026 32564
rect 617 32527 1026 32530
rect 617 32496 814 32527
rect 617 32462 646 32496
rect 680 32493 814 32496
rect 848 32493 1026 32527
rect 680 32462 1026 32493
rect 617 32455 1026 32462
rect 617 32428 814 32455
rect 617 32394 646 32428
rect 680 32421 814 32428
rect 848 32421 1026 32455
rect 680 32394 1026 32421
rect 617 32383 1026 32394
rect 617 32360 814 32383
rect 617 32326 646 32360
rect 680 32349 814 32360
rect 848 32349 1026 32383
rect 680 32326 1026 32349
rect 617 32311 1026 32326
rect 617 32292 814 32311
rect 617 32258 646 32292
rect 680 32277 814 32292
rect 848 32277 1026 32311
rect 680 32258 1026 32277
rect 617 32239 1026 32258
rect 617 32224 814 32239
rect 617 32190 646 32224
rect 680 32205 814 32224
rect 848 32205 1026 32239
rect 680 32190 1026 32205
rect 617 32167 1026 32190
rect 617 32156 814 32167
rect 617 32122 646 32156
rect 680 32133 814 32156
rect 848 32133 1026 32167
rect 680 32122 1026 32133
rect 617 32095 1026 32122
rect 617 32088 814 32095
rect 617 32054 646 32088
rect 680 32061 814 32088
rect 848 32061 1026 32095
rect 680 32054 1026 32061
rect 617 32023 1026 32054
rect 617 32020 814 32023
rect 617 31986 646 32020
rect 680 31989 814 32020
rect 848 31989 1026 32023
rect 680 31986 1026 31989
rect 617 31952 1026 31986
rect 617 31918 646 31952
rect 680 31951 1026 31952
rect 680 31918 814 31951
rect 617 31917 814 31918
rect 848 31917 1026 31951
rect 617 31884 1026 31917
rect 617 31850 646 31884
rect 680 31879 1026 31884
rect 680 31850 814 31879
rect 617 31845 814 31850
rect 848 31845 1026 31879
rect 617 31816 1026 31845
rect 617 31782 646 31816
rect 680 31807 1026 31816
rect 680 31782 814 31807
rect 617 31773 814 31782
rect 848 31773 1026 31807
rect 617 31748 1026 31773
rect 617 31714 646 31748
rect 680 31735 1026 31748
rect 680 31714 814 31735
rect 617 31701 814 31714
rect 848 31701 1026 31735
rect 617 31680 1026 31701
rect 617 31646 646 31680
rect 680 31663 1026 31680
rect 680 31646 814 31663
rect 617 31629 814 31646
rect 848 31629 1026 31663
rect 617 31612 1026 31629
rect 617 31578 646 31612
rect 680 31591 1026 31612
rect 680 31578 814 31591
rect 617 31557 814 31578
rect 848 31557 1026 31591
rect 617 31544 1026 31557
rect 617 31510 646 31544
rect 680 31519 1026 31544
rect 680 31510 814 31519
rect 617 31485 814 31510
rect 848 31485 1026 31519
rect 617 31476 1026 31485
rect 617 31442 646 31476
rect 680 31447 1026 31476
rect 680 31442 814 31447
rect 617 31413 814 31442
rect 848 31413 1026 31447
rect 617 31408 1026 31413
rect 617 31374 646 31408
rect 680 31375 1026 31408
rect 680 31374 814 31375
rect 617 31341 814 31374
rect 848 31341 1026 31375
rect 617 31340 1026 31341
rect 617 31306 646 31340
rect 680 31306 1026 31340
rect 617 31303 1026 31306
rect 617 31272 814 31303
rect 617 31238 646 31272
rect 680 31269 814 31272
rect 848 31269 1026 31303
rect 680 31238 1026 31269
rect 617 31231 1026 31238
rect 617 31204 814 31231
rect 617 31170 646 31204
rect 680 31197 814 31204
rect 848 31197 1026 31231
rect 680 31170 1026 31197
rect 617 31159 1026 31170
rect 617 31136 814 31159
rect 617 31102 646 31136
rect 680 31125 814 31136
rect 848 31125 1026 31159
rect 680 31102 1026 31125
rect 617 31087 1026 31102
rect 617 31068 814 31087
rect 617 31034 646 31068
rect 680 31053 814 31068
rect 848 31053 1026 31087
rect 680 31034 1026 31053
rect 617 31015 1026 31034
rect 617 31000 814 31015
rect 617 30966 646 31000
rect 680 30981 814 31000
rect 848 30981 1026 31015
rect 680 30966 1026 30981
rect 617 30943 1026 30966
rect 617 30932 814 30943
rect 617 30898 646 30932
rect 680 30909 814 30932
rect 848 30909 1026 30943
rect 680 30898 1026 30909
rect 617 30871 1026 30898
rect 617 30864 814 30871
rect 617 30830 646 30864
rect 680 30837 814 30864
rect 848 30837 1026 30871
rect 680 30830 1026 30837
rect 617 30799 1026 30830
rect 617 30796 814 30799
rect 617 30762 646 30796
rect 680 30765 814 30796
rect 848 30765 1026 30799
rect 680 30762 1026 30765
rect 617 30728 1026 30762
rect 617 30694 646 30728
rect 680 30727 1026 30728
rect 680 30694 814 30727
rect 617 30693 814 30694
rect 848 30693 1026 30727
rect 617 30660 1026 30693
rect 617 30626 646 30660
rect 680 30655 1026 30660
rect 680 30626 814 30655
rect 617 30621 814 30626
rect 848 30621 1026 30655
rect 617 30592 1026 30621
rect 617 30558 646 30592
rect 680 30583 1026 30592
rect 680 30558 814 30583
rect 617 30549 814 30558
rect 848 30549 1026 30583
rect 617 30524 1026 30549
rect 617 30490 646 30524
rect 680 30511 1026 30524
rect 680 30490 814 30511
rect 617 30477 814 30490
rect 848 30477 1026 30511
rect 617 30456 1026 30477
rect 617 30422 646 30456
rect 680 30439 1026 30456
rect 680 30422 814 30439
rect 617 30405 814 30422
rect 848 30405 1026 30439
rect 617 30388 1026 30405
rect 617 30354 646 30388
rect 680 30367 1026 30388
rect 680 30354 814 30367
rect 617 30333 814 30354
rect 848 30333 1026 30367
rect 617 30320 1026 30333
rect 617 30286 646 30320
rect 680 30295 1026 30320
rect 680 30286 814 30295
rect 617 30261 814 30286
rect 848 30261 1026 30295
rect 617 30252 1026 30261
rect 617 30218 646 30252
rect 680 30223 1026 30252
rect 680 30218 814 30223
rect 617 30189 814 30218
rect 848 30189 1026 30223
rect 617 30184 1026 30189
rect 617 30150 646 30184
rect 680 30151 1026 30184
rect 680 30150 814 30151
rect 617 30117 814 30150
rect 848 30117 1026 30151
rect 617 30116 1026 30117
rect 617 30082 646 30116
rect 680 30082 1026 30116
rect 617 30079 1026 30082
rect 617 30048 814 30079
rect 617 30014 646 30048
rect 680 30045 814 30048
rect 848 30045 1026 30079
rect 680 30014 1026 30045
rect 617 30007 1026 30014
rect 617 29980 814 30007
rect 617 29946 646 29980
rect 680 29973 814 29980
rect 848 29973 1026 30007
rect 680 29946 1026 29973
rect 617 29935 1026 29946
rect 617 29912 814 29935
rect 617 29878 646 29912
rect 680 29901 814 29912
rect 848 29901 1026 29935
rect 680 29878 1026 29901
rect 617 29863 1026 29878
rect 617 29844 814 29863
rect 617 29810 646 29844
rect 680 29829 814 29844
rect 848 29829 1026 29863
rect 680 29810 1026 29829
rect 617 29791 1026 29810
rect 617 29776 814 29791
rect 617 29742 646 29776
rect 680 29757 814 29776
rect 848 29757 1026 29791
rect 680 29742 1026 29757
rect 617 29719 1026 29742
rect 617 29708 814 29719
rect 617 29674 646 29708
rect 680 29685 814 29708
rect 848 29685 1026 29719
rect 680 29674 1026 29685
rect 617 29647 1026 29674
rect 617 29640 814 29647
rect 617 29606 646 29640
rect 680 29613 814 29640
rect 848 29613 1026 29647
rect 680 29606 1026 29613
rect 617 29575 1026 29606
rect 617 29572 814 29575
rect 617 29538 646 29572
rect 680 29541 814 29572
rect 848 29541 1026 29575
rect 680 29538 1026 29541
rect 617 29504 1026 29538
rect 617 29470 646 29504
rect 680 29503 1026 29504
rect 680 29470 814 29503
rect 617 29469 814 29470
rect 848 29469 1026 29503
rect 617 29436 1026 29469
rect 617 29402 646 29436
rect 680 29431 1026 29436
rect 680 29402 814 29431
rect 617 29397 814 29402
rect 848 29397 1026 29431
rect 617 29368 1026 29397
rect 617 29334 646 29368
rect 680 29359 1026 29368
rect 680 29334 814 29359
rect 617 29325 814 29334
rect 848 29325 1026 29359
rect 617 29300 1026 29325
rect 617 29266 646 29300
rect 680 29287 1026 29300
rect 680 29266 814 29287
rect 617 29253 814 29266
rect 848 29253 1026 29287
rect 617 29232 1026 29253
rect 617 29198 646 29232
rect 680 29215 1026 29232
rect 680 29198 814 29215
rect 617 29181 814 29198
rect 848 29181 1026 29215
rect 617 29164 1026 29181
rect 617 29130 646 29164
rect 680 29143 1026 29164
rect 680 29130 814 29143
rect 617 29109 814 29130
rect 848 29109 1026 29143
rect 617 29096 1026 29109
rect 617 29062 646 29096
rect 680 29071 1026 29096
rect 680 29062 814 29071
rect 617 29037 814 29062
rect 848 29037 1026 29071
rect 617 29028 1026 29037
rect 617 28994 646 29028
rect 680 28999 1026 29028
rect 680 28994 814 28999
rect 617 28965 814 28994
rect 848 28965 1026 28999
rect 617 28960 1026 28965
rect 617 28926 646 28960
rect 680 28927 1026 28960
rect 680 28926 814 28927
rect 617 28893 814 28926
rect 848 28893 1026 28927
rect 617 28892 1026 28893
rect 617 28858 646 28892
rect 680 28858 1026 28892
rect 617 28855 1026 28858
rect 617 28824 814 28855
rect 617 28790 646 28824
rect 680 28821 814 28824
rect 848 28821 1026 28855
rect 680 28790 1026 28821
rect 617 28783 1026 28790
rect 617 28756 814 28783
rect 617 28722 646 28756
rect 680 28749 814 28756
rect 848 28749 1026 28783
rect 680 28722 1026 28749
rect 617 28711 1026 28722
rect 617 28688 814 28711
rect 617 28654 646 28688
rect 680 28677 814 28688
rect 848 28677 1026 28711
rect 680 28654 1026 28677
rect 617 28639 1026 28654
rect 617 28620 814 28639
rect 617 28586 646 28620
rect 680 28605 814 28620
rect 848 28605 1026 28639
rect 680 28586 1026 28605
rect 617 28567 1026 28586
rect 617 28552 814 28567
rect 617 28518 646 28552
rect 680 28533 814 28552
rect 848 28533 1026 28567
rect 680 28518 1026 28533
rect 617 28495 1026 28518
rect 617 28484 814 28495
rect 617 28450 646 28484
rect 680 28461 814 28484
rect 848 28461 1026 28495
rect 680 28450 1026 28461
rect 617 28423 1026 28450
rect 617 28416 814 28423
rect 617 28382 646 28416
rect 680 28389 814 28416
rect 848 28389 1026 28423
rect 680 28382 1026 28389
rect 617 28351 1026 28382
rect 617 28348 814 28351
rect 617 28314 646 28348
rect 680 28317 814 28348
rect 848 28317 1026 28351
rect 680 28314 1026 28317
rect 617 28280 1026 28314
rect 617 28246 646 28280
rect 680 28279 1026 28280
rect 680 28246 814 28279
rect 617 28245 814 28246
rect 848 28245 1026 28279
rect 617 28212 1026 28245
rect 617 28178 646 28212
rect 680 28207 1026 28212
rect 680 28178 814 28207
rect 617 28173 814 28178
rect 848 28173 1026 28207
rect 617 28144 1026 28173
rect 617 28110 646 28144
rect 680 28135 1026 28144
rect 680 28110 814 28135
rect 617 28101 814 28110
rect 848 28101 1026 28135
rect 617 28076 1026 28101
rect 617 28042 646 28076
rect 680 28063 1026 28076
rect 680 28042 814 28063
rect 617 28029 814 28042
rect 848 28029 1026 28063
rect 617 28008 1026 28029
rect 617 27974 646 28008
rect 680 27991 1026 28008
rect 680 27974 814 27991
rect 617 27957 814 27974
rect 848 27957 1026 27991
rect 617 27940 1026 27957
rect 617 27906 646 27940
rect 680 27919 1026 27940
rect 680 27906 814 27919
rect 617 27885 814 27906
rect 848 27885 1026 27919
rect 617 27872 1026 27885
rect 617 27838 646 27872
rect 680 27847 1026 27872
rect 680 27838 814 27847
rect 617 27813 814 27838
rect 848 27813 1026 27847
rect 617 27804 1026 27813
rect 617 27770 646 27804
rect 680 27775 1026 27804
rect 680 27770 814 27775
rect 617 27741 814 27770
rect 848 27741 1026 27775
rect 617 27736 1026 27741
rect 617 27702 646 27736
rect 680 27703 1026 27736
rect 680 27702 814 27703
rect 617 27669 814 27702
rect 848 27669 1026 27703
rect 617 27668 1026 27669
rect 617 27634 646 27668
rect 680 27634 1026 27668
rect 617 27631 1026 27634
rect 617 27600 814 27631
rect 617 27566 646 27600
rect 680 27597 814 27600
rect 848 27597 1026 27631
rect 680 27566 1026 27597
rect 617 27559 1026 27566
rect 617 27532 814 27559
rect 617 27498 646 27532
rect 680 27525 814 27532
rect 848 27525 1026 27559
rect 680 27498 1026 27525
rect 617 27487 1026 27498
rect 617 27464 814 27487
rect 617 27430 646 27464
rect 680 27453 814 27464
rect 848 27453 1026 27487
rect 680 27430 1026 27453
rect 617 27415 1026 27430
rect 617 27396 814 27415
rect 617 27362 646 27396
rect 680 27381 814 27396
rect 848 27381 1026 27415
rect 680 27362 1026 27381
rect 617 27343 1026 27362
rect 617 27328 814 27343
rect 617 27294 646 27328
rect 680 27309 814 27328
rect 848 27309 1026 27343
rect 680 27294 1026 27309
rect 617 27271 1026 27294
rect 617 27260 814 27271
rect 617 27226 646 27260
rect 680 27237 814 27260
rect 848 27237 1026 27271
rect 680 27226 1026 27237
rect 617 27199 1026 27226
rect 617 27192 814 27199
rect 617 27158 646 27192
rect 680 27165 814 27192
rect 848 27165 1026 27199
rect 680 27158 1026 27165
rect 617 27127 1026 27158
rect 617 27124 814 27127
rect 617 27090 646 27124
rect 680 27093 814 27124
rect 848 27093 1026 27127
rect 680 27090 1026 27093
rect 617 27056 1026 27090
rect 617 27022 646 27056
rect 680 27055 1026 27056
rect 680 27022 814 27055
rect 617 27021 814 27022
rect 848 27021 1026 27055
rect 617 26988 1026 27021
rect 617 26954 646 26988
rect 680 26983 1026 26988
rect 680 26954 814 26983
rect 617 26949 814 26954
rect 848 26949 1026 26983
rect 617 26920 1026 26949
rect 617 26886 646 26920
rect 680 26911 1026 26920
rect 680 26886 814 26911
rect 617 26877 814 26886
rect 848 26877 1026 26911
rect 617 26852 1026 26877
rect 617 26818 646 26852
rect 680 26839 1026 26852
rect 680 26818 814 26839
rect 617 26805 814 26818
rect 848 26805 1026 26839
rect 617 26784 1026 26805
rect 617 26750 646 26784
rect 680 26767 1026 26784
rect 680 26750 814 26767
rect 617 26733 814 26750
rect 848 26733 1026 26767
rect 617 26716 1026 26733
rect 617 26682 646 26716
rect 680 26695 1026 26716
rect 680 26682 814 26695
rect 617 26661 814 26682
rect 848 26661 1026 26695
rect 617 26648 1026 26661
rect 617 26614 646 26648
rect 680 26623 1026 26648
rect 680 26614 814 26623
rect 617 26589 814 26614
rect 848 26589 1026 26623
rect 617 26580 1026 26589
rect 617 26546 646 26580
rect 680 26551 1026 26580
rect 680 26546 814 26551
rect 617 26517 814 26546
rect 848 26517 1026 26551
rect 617 26512 1026 26517
rect 617 26478 646 26512
rect 680 26479 1026 26512
rect 680 26478 814 26479
rect 617 26445 814 26478
rect 848 26445 1026 26479
rect 617 26444 1026 26445
rect 617 26410 646 26444
rect 680 26410 1026 26444
rect 617 26407 1026 26410
rect 617 26376 814 26407
rect 617 26342 646 26376
rect 680 26373 814 26376
rect 848 26373 1026 26407
rect 680 26342 1026 26373
rect 617 26335 1026 26342
rect 617 26308 814 26335
rect 617 26274 646 26308
rect 680 26301 814 26308
rect 848 26301 1026 26335
rect 680 26274 1026 26301
rect 617 26263 1026 26274
rect 617 26240 814 26263
rect 617 26206 646 26240
rect 680 26229 814 26240
rect 848 26229 1026 26263
rect 680 26206 1026 26229
rect 617 26191 1026 26206
rect 617 26172 814 26191
rect 617 26138 646 26172
rect 680 26157 814 26172
rect 848 26157 1026 26191
rect 680 26138 1026 26157
rect 617 26119 1026 26138
rect 617 26104 814 26119
rect 617 26070 646 26104
rect 680 26085 814 26104
rect 848 26085 1026 26119
rect 680 26070 1026 26085
rect 617 26047 1026 26070
rect 617 26036 814 26047
rect 617 26002 646 26036
rect 680 26013 814 26036
rect 848 26013 1026 26047
rect 680 26002 1026 26013
rect 617 25975 1026 26002
rect 617 25968 814 25975
rect 617 25934 646 25968
rect 680 25941 814 25968
rect 848 25941 1026 25975
rect 680 25934 1026 25941
rect 617 25903 1026 25934
rect 617 25900 814 25903
rect 617 25866 646 25900
rect 680 25869 814 25900
rect 848 25869 1026 25903
rect 680 25866 1026 25869
rect 617 25832 1026 25866
rect 617 25798 646 25832
rect 680 25831 1026 25832
rect 680 25798 814 25831
rect 617 25797 814 25798
rect 848 25797 1026 25831
rect 617 25764 1026 25797
rect 617 25730 646 25764
rect 680 25759 1026 25764
rect 680 25730 814 25759
rect 617 25725 814 25730
rect 848 25725 1026 25759
rect 617 25696 1026 25725
rect 617 25662 646 25696
rect 680 25687 1026 25696
rect 680 25662 814 25687
rect 617 25653 814 25662
rect 848 25653 1026 25687
rect 617 25628 1026 25653
rect 617 25594 646 25628
rect 680 25615 1026 25628
rect 680 25594 814 25615
rect 617 25581 814 25594
rect 848 25581 1026 25615
rect 617 25560 1026 25581
rect 617 25526 646 25560
rect 680 25543 1026 25560
rect 680 25526 814 25543
rect 617 25509 814 25526
rect 848 25509 1026 25543
rect 617 25492 1026 25509
rect 617 25458 646 25492
rect 680 25471 1026 25492
rect 680 25458 814 25471
rect 617 25437 814 25458
rect 848 25437 1026 25471
rect 617 25424 1026 25437
rect 617 25390 646 25424
rect 680 25399 1026 25424
rect 680 25390 814 25399
rect 617 25365 814 25390
rect 848 25365 1026 25399
rect 617 25356 1026 25365
rect 617 25322 646 25356
rect 680 25327 1026 25356
rect 680 25322 814 25327
rect 617 25293 814 25322
rect 848 25293 1026 25327
rect 617 25288 1026 25293
rect 617 25254 646 25288
rect 680 25255 1026 25288
rect 680 25254 814 25255
rect 617 25221 814 25254
rect 848 25221 1026 25255
rect 617 25220 1026 25221
rect 617 25186 646 25220
rect 680 25186 1026 25220
rect 617 25183 1026 25186
rect 617 25152 814 25183
rect 617 25118 646 25152
rect 680 25149 814 25152
rect 848 25149 1026 25183
rect 680 25118 1026 25149
rect 617 25111 1026 25118
rect 617 25084 814 25111
rect 617 25050 646 25084
rect 680 25077 814 25084
rect 848 25077 1026 25111
rect 680 25050 1026 25077
rect 617 25039 1026 25050
rect 617 25016 814 25039
rect 617 24982 646 25016
rect 680 25005 814 25016
rect 848 25005 1026 25039
rect 680 24982 1026 25005
rect 617 24967 1026 24982
rect 617 24948 814 24967
rect 617 24914 646 24948
rect 680 24933 814 24948
rect 848 24933 1026 24967
rect 680 24914 1026 24933
rect 617 24895 1026 24914
rect 617 24880 814 24895
rect 617 24846 646 24880
rect 680 24861 814 24880
rect 848 24861 1026 24895
rect 680 24846 1026 24861
rect 617 24823 1026 24846
rect 617 24812 814 24823
rect 617 24778 646 24812
rect 680 24789 814 24812
rect 848 24789 1026 24823
rect 680 24778 1026 24789
rect 617 24751 1026 24778
rect 617 24744 814 24751
rect 617 24710 646 24744
rect 680 24717 814 24744
rect 848 24717 1026 24751
rect 680 24710 1026 24717
rect 617 24679 1026 24710
rect 617 24676 814 24679
rect 617 24642 646 24676
rect 680 24645 814 24676
rect 848 24645 1026 24679
rect 680 24642 1026 24645
rect 617 24608 1026 24642
rect 617 24574 646 24608
rect 680 24607 1026 24608
rect 680 24574 814 24607
rect 617 24573 814 24574
rect 848 24573 1026 24607
rect 617 24540 1026 24573
rect 617 24506 646 24540
rect 680 24535 1026 24540
rect 680 24506 814 24535
rect 617 24501 814 24506
rect 848 24501 1026 24535
rect 617 24472 1026 24501
rect 617 24438 646 24472
rect 680 24463 1026 24472
rect 680 24438 814 24463
rect 617 24429 814 24438
rect 848 24429 1026 24463
rect 617 24404 1026 24429
rect 617 24370 646 24404
rect 680 24391 1026 24404
rect 680 24370 814 24391
rect 617 24357 814 24370
rect 848 24357 1026 24391
rect 617 24336 1026 24357
rect 617 24302 646 24336
rect 680 24319 1026 24336
rect 680 24302 814 24319
rect 617 24285 814 24302
rect 848 24285 1026 24319
rect 617 24268 1026 24285
rect 617 24234 646 24268
rect 680 24247 1026 24268
rect 680 24234 814 24247
rect 617 24213 814 24234
rect 848 24213 1026 24247
rect 617 24200 1026 24213
rect 617 24166 646 24200
rect 680 24175 1026 24200
rect 680 24166 814 24175
rect 617 24141 814 24166
rect 848 24141 1026 24175
rect 617 24132 1026 24141
rect 617 24098 646 24132
rect 680 24103 1026 24132
rect 680 24098 814 24103
rect 617 24069 814 24098
rect 848 24069 1026 24103
rect 617 24064 1026 24069
rect 617 24030 646 24064
rect 680 24031 1026 24064
rect 680 24030 814 24031
rect 617 23997 814 24030
rect 848 23997 1026 24031
rect 617 23996 1026 23997
rect 617 23962 646 23996
rect 680 23962 1026 23996
rect 617 23959 1026 23962
rect 617 23928 814 23959
rect 617 23894 646 23928
rect 680 23925 814 23928
rect 848 23925 1026 23959
rect 680 23894 1026 23925
rect 617 23887 1026 23894
rect 617 23860 814 23887
rect 617 23826 646 23860
rect 680 23853 814 23860
rect 848 23853 1026 23887
rect 680 23826 1026 23853
rect 617 23815 1026 23826
rect 617 23792 814 23815
rect 617 23758 646 23792
rect 680 23781 814 23792
rect 848 23781 1026 23815
rect 680 23758 1026 23781
rect 617 23743 1026 23758
rect 617 23724 814 23743
rect 617 23690 646 23724
rect 680 23709 814 23724
rect 848 23709 1026 23743
rect 680 23690 1026 23709
rect 617 23671 1026 23690
rect 617 23656 814 23671
rect 617 23622 646 23656
rect 680 23637 814 23656
rect 848 23637 1026 23671
rect 680 23622 1026 23637
rect 617 23599 1026 23622
rect 617 23588 814 23599
rect 617 23554 646 23588
rect 680 23565 814 23588
rect 848 23565 1026 23599
rect 680 23554 1026 23565
rect 617 23527 1026 23554
rect 617 23520 814 23527
rect 617 23486 646 23520
rect 680 23493 814 23520
rect 848 23493 1026 23527
rect 680 23486 1026 23493
rect 617 23455 1026 23486
rect 617 23452 814 23455
rect 617 23418 646 23452
rect 680 23421 814 23452
rect 848 23421 1026 23455
rect 680 23418 1026 23421
rect 617 23384 1026 23418
rect 617 23350 646 23384
rect 680 23383 1026 23384
rect 680 23350 814 23383
rect 617 23349 814 23350
rect 848 23349 1026 23383
rect 617 23316 1026 23349
rect 617 23282 646 23316
rect 680 23311 1026 23316
rect 680 23282 814 23311
rect 617 23277 814 23282
rect 848 23277 1026 23311
rect 617 23248 1026 23277
rect 617 23214 646 23248
rect 680 23239 1026 23248
rect 680 23214 814 23239
rect 617 23205 814 23214
rect 848 23205 1026 23239
rect 617 23180 1026 23205
rect 617 23146 646 23180
rect 680 23167 1026 23180
rect 680 23146 814 23167
rect 617 23133 814 23146
rect 848 23133 1026 23167
rect 617 23112 1026 23133
rect 617 23078 646 23112
rect 680 23095 1026 23112
rect 680 23078 814 23095
rect 617 23061 814 23078
rect 848 23061 1026 23095
rect 617 23044 1026 23061
rect 617 23010 646 23044
rect 680 23023 1026 23044
rect 680 23010 814 23023
rect 617 22989 814 23010
rect 848 22989 1026 23023
rect 617 22976 1026 22989
rect 617 22942 646 22976
rect 680 22951 1026 22976
rect 680 22942 814 22951
rect 617 22917 814 22942
rect 848 22917 1026 22951
rect 617 22908 1026 22917
rect 617 22874 646 22908
rect 680 22879 1026 22908
rect 680 22874 814 22879
rect 617 22845 814 22874
rect 848 22845 1026 22879
rect 617 22840 1026 22845
rect 617 22806 646 22840
rect 680 22807 1026 22840
rect 680 22806 814 22807
rect 617 22773 814 22806
rect 848 22773 1026 22807
rect 617 22772 1026 22773
rect 617 22738 646 22772
rect 680 22738 1026 22772
rect 617 22735 1026 22738
rect 617 22704 814 22735
rect 617 22670 646 22704
rect 680 22701 814 22704
rect 848 22701 1026 22735
rect 680 22670 1026 22701
rect 617 22663 1026 22670
rect 617 22636 814 22663
rect 617 22602 646 22636
rect 680 22629 814 22636
rect 848 22629 1026 22663
rect 680 22602 1026 22629
rect 617 22591 1026 22602
rect 617 22568 814 22591
rect 617 22534 646 22568
rect 680 22557 814 22568
rect 848 22557 1026 22591
rect 680 22534 1026 22557
rect 617 22519 1026 22534
rect 617 22500 814 22519
rect 617 22466 646 22500
rect 680 22485 814 22500
rect 848 22485 1026 22519
rect 680 22466 1026 22485
rect 617 22447 1026 22466
rect 617 22432 814 22447
rect 617 22398 646 22432
rect 680 22413 814 22432
rect 848 22413 1026 22447
rect 680 22398 1026 22413
rect 617 22375 1026 22398
rect 617 22364 814 22375
rect 617 22330 646 22364
rect 680 22341 814 22364
rect 848 22341 1026 22375
rect 680 22330 1026 22341
rect 617 22303 1026 22330
rect 617 22296 814 22303
rect 617 22262 646 22296
rect 680 22269 814 22296
rect 848 22269 1026 22303
rect 680 22262 1026 22269
rect 617 22231 1026 22262
rect 617 22228 814 22231
rect 617 22194 646 22228
rect 680 22197 814 22228
rect 848 22197 1026 22231
rect 680 22194 1026 22197
rect 617 22160 1026 22194
rect 617 22126 646 22160
rect 680 22159 1026 22160
rect 680 22126 814 22159
rect 617 22125 814 22126
rect 848 22125 1026 22159
rect 617 22092 1026 22125
rect 617 22058 646 22092
rect 680 22087 1026 22092
rect 680 22058 814 22087
rect 617 22053 814 22058
rect 848 22053 1026 22087
rect 617 22024 1026 22053
rect 617 21990 646 22024
rect 680 22015 1026 22024
rect 680 21990 814 22015
rect 617 21981 814 21990
rect 848 21981 1026 22015
rect 617 21956 1026 21981
rect 617 21922 646 21956
rect 680 21943 1026 21956
rect 680 21922 814 21943
rect 617 21909 814 21922
rect 848 21909 1026 21943
rect 617 21888 1026 21909
rect 617 21854 646 21888
rect 680 21871 1026 21888
rect 680 21854 814 21871
rect 617 21837 814 21854
rect 848 21837 1026 21871
rect 617 21820 1026 21837
rect 617 21786 646 21820
rect 680 21799 1026 21820
rect 680 21786 814 21799
rect 617 21765 814 21786
rect 848 21765 1026 21799
rect 617 21752 1026 21765
rect 617 21718 646 21752
rect 680 21727 1026 21752
rect 680 21718 814 21727
rect 617 21693 814 21718
rect 848 21693 1026 21727
rect 617 21684 1026 21693
rect 617 21650 646 21684
rect 680 21655 1026 21684
rect 680 21650 814 21655
rect 617 21621 814 21650
rect 848 21621 1026 21655
rect 617 21616 1026 21621
rect 617 21582 646 21616
rect 680 21583 1026 21616
rect 680 21582 814 21583
rect 617 21549 814 21582
rect 848 21549 1026 21583
rect 617 21548 1026 21549
rect 617 21514 646 21548
rect 680 21514 1026 21548
rect 617 21511 1026 21514
rect 617 21480 814 21511
rect 617 21446 646 21480
rect 680 21477 814 21480
rect 848 21477 1026 21511
rect 680 21446 1026 21477
rect 617 21439 1026 21446
rect 617 21412 814 21439
rect 617 21378 646 21412
rect 680 21405 814 21412
rect 848 21405 1026 21439
rect 680 21378 1026 21405
rect 617 21367 1026 21378
rect 617 21344 814 21367
rect 617 21310 646 21344
rect 680 21333 814 21344
rect 848 21333 1026 21367
rect 680 21310 1026 21333
rect 617 21295 1026 21310
rect 617 21276 814 21295
rect 617 21242 646 21276
rect 680 21261 814 21276
rect 848 21261 1026 21295
rect 680 21242 1026 21261
rect 617 21223 1026 21242
rect 617 21208 814 21223
rect 617 21174 646 21208
rect 680 21189 814 21208
rect 848 21189 1026 21223
rect 680 21174 1026 21189
rect 617 21151 1026 21174
rect 617 21140 814 21151
rect 617 21106 646 21140
rect 680 21117 814 21140
rect 848 21117 1026 21151
rect 680 21106 1026 21117
rect 617 21079 1026 21106
rect 617 21072 814 21079
rect 617 21038 646 21072
rect 680 21045 814 21072
rect 848 21045 1026 21079
rect 680 21038 1026 21045
rect 617 21007 1026 21038
rect 617 21004 814 21007
rect 617 20970 646 21004
rect 680 20973 814 21004
rect 848 20973 1026 21007
rect 680 20970 1026 20973
rect 617 20936 1026 20970
rect 617 20902 646 20936
rect 680 20935 1026 20936
rect 680 20902 814 20935
rect 617 20901 814 20902
rect 848 20901 1026 20935
rect 617 20868 1026 20901
rect 617 20834 646 20868
rect 680 20863 1026 20868
rect 680 20834 814 20863
rect 617 20829 814 20834
rect 848 20829 1026 20863
rect 617 20800 1026 20829
rect 617 20766 646 20800
rect 680 20791 1026 20800
rect 680 20766 814 20791
rect 617 20757 814 20766
rect 848 20757 1026 20791
rect 617 20732 1026 20757
rect 617 20698 646 20732
rect 680 20719 1026 20732
rect 680 20698 814 20719
rect 617 20685 814 20698
rect 848 20685 1026 20719
rect 617 20664 1026 20685
rect 617 20630 646 20664
rect 680 20647 1026 20664
rect 680 20630 814 20647
rect 617 20613 814 20630
rect 848 20613 1026 20647
rect 617 20596 1026 20613
rect 617 20562 646 20596
rect 680 20575 1026 20596
rect 680 20562 814 20575
rect 617 20541 814 20562
rect 848 20541 1026 20575
rect 617 20528 1026 20541
rect 617 20494 646 20528
rect 680 20503 1026 20528
rect 680 20494 814 20503
rect 617 20469 814 20494
rect 848 20469 1026 20503
rect 617 20460 1026 20469
rect 617 20426 646 20460
rect 680 20431 1026 20460
rect 680 20426 814 20431
rect 617 20397 814 20426
rect 848 20397 1026 20431
rect 617 20392 1026 20397
rect 617 20358 646 20392
rect 680 20359 1026 20392
rect 680 20358 814 20359
rect 617 20325 814 20358
rect 848 20325 1026 20359
rect 617 20324 1026 20325
rect 617 20290 646 20324
rect 680 20290 1026 20324
rect 617 20287 1026 20290
rect 617 20256 814 20287
rect 617 20222 646 20256
rect 680 20253 814 20256
rect 848 20253 1026 20287
rect 680 20222 1026 20253
rect 617 20215 1026 20222
rect 617 20188 814 20215
rect 617 20154 646 20188
rect 680 20181 814 20188
rect 848 20181 1026 20215
rect 680 20154 1026 20181
rect 617 20143 1026 20154
rect 617 20120 814 20143
rect 617 20086 646 20120
rect 680 20109 814 20120
rect 848 20109 1026 20143
rect 680 20086 1026 20109
rect 617 20071 1026 20086
rect 617 20052 814 20071
rect 617 20018 646 20052
rect 680 20037 814 20052
rect 848 20037 1026 20071
rect 680 20018 1026 20037
rect 617 19999 1026 20018
rect 617 19984 814 19999
rect 617 19950 646 19984
rect 680 19965 814 19984
rect 848 19965 1026 19999
rect 680 19950 1026 19965
rect 617 19927 1026 19950
rect 617 19916 814 19927
rect 617 19882 646 19916
rect 680 19893 814 19916
rect 848 19893 1026 19927
rect 680 19882 1026 19893
rect 617 19855 1026 19882
rect 617 19848 814 19855
rect 617 19814 646 19848
rect 680 19821 814 19848
rect 848 19821 1026 19855
rect 680 19814 1026 19821
rect 617 19783 1026 19814
rect 617 19780 814 19783
rect 617 19746 646 19780
rect 680 19749 814 19780
rect 848 19749 1026 19783
rect 680 19746 1026 19749
rect 617 19712 1026 19746
rect 617 19678 646 19712
rect 680 19711 1026 19712
rect 680 19678 814 19711
rect 617 19677 814 19678
rect 848 19677 1026 19711
rect 617 19644 1026 19677
rect 617 19610 646 19644
rect 680 19639 1026 19644
rect 680 19610 814 19639
rect 617 19605 814 19610
rect 848 19605 1026 19639
rect 617 19576 1026 19605
rect 617 19542 646 19576
rect 680 19567 1026 19576
rect 680 19542 814 19567
rect 617 19533 814 19542
rect 848 19533 1026 19567
rect 617 19508 1026 19533
rect 617 19474 646 19508
rect 680 19495 1026 19508
rect 680 19474 814 19495
rect 617 19461 814 19474
rect 848 19461 1026 19495
rect 617 19440 1026 19461
rect 617 19406 646 19440
rect 680 19423 1026 19440
rect 680 19406 814 19423
rect 617 19389 814 19406
rect 848 19389 1026 19423
rect 617 19372 1026 19389
rect 617 19338 646 19372
rect 680 19351 1026 19372
rect 680 19338 814 19351
rect 617 19317 814 19338
rect 848 19317 1026 19351
rect 617 19304 1026 19317
rect 617 19270 646 19304
rect 680 19279 1026 19304
rect 680 19270 814 19279
rect 617 19245 814 19270
rect 848 19245 1026 19279
rect 617 19236 1026 19245
rect 617 19202 646 19236
rect 680 19207 1026 19236
rect 680 19202 814 19207
rect 617 19173 814 19202
rect 848 19173 1026 19207
rect 617 19168 1026 19173
rect 617 19134 646 19168
rect 680 19135 1026 19168
rect 680 19134 814 19135
rect 617 19101 814 19134
rect 848 19101 1026 19135
rect 617 19100 1026 19101
rect 617 19066 646 19100
rect 680 19066 1026 19100
rect 617 19063 1026 19066
rect 617 19032 814 19063
rect 617 18998 646 19032
rect 680 19029 814 19032
rect 848 19029 1026 19063
rect 680 18998 1026 19029
rect 617 18991 1026 18998
rect 617 18964 814 18991
rect 617 18930 646 18964
rect 680 18957 814 18964
rect 848 18957 1026 18991
rect 680 18930 1026 18957
rect 617 18919 1026 18930
rect 617 18896 814 18919
rect 617 18862 646 18896
rect 680 18885 814 18896
rect 848 18885 1026 18919
rect 680 18862 1026 18885
rect 617 18847 1026 18862
rect 617 18828 814 18847
rect 617 18794 646 18828
rect 680 18813 814 18828
rect 848 18813 1026 18847
rect 680 18794 1026 18813
rect 617 18775 1026 18794
rect 617 18760 814 18775
rect 617 18726 646 18760
rect 680 18741 814 18760
rect 848 18741 1026 18775
rect 680 18726 1026 18741
rect 617 18703 1026 18726
rect 617 18692 814 18703
rect 617 18658 646 18692
rect 680 18669 814 18692
rect 848 18669 1026 18703
rect 680 18658 1026 18669
rect 617 18631 1026 18658
rect 617 18624 814 18631
rect 617 18590 646 18624
rect 680 18597 814 18624
rect 848 18597 1026 18631
rect 680 18590 1026 18597
rect 617 18559 1026 18590
rect 617 18556 814 18559
rect 617 18522 646 18556
rect 680 18525 814 18556
rect 848 18525 1026 18559
rect 680 18522 1026 18525
rect 617 18488 1026 18522
rect 617 18454 646 18488
rect 680 18487 1026 18488
rect 680 18454 814 18487
rect 617 18453 814 18454
rect 848 18453 1026 18487
rect 617 18420 1026 18453
rect 617 18386 646 18420
rect 680 18415 1026 18420
rect 680 18386 814 18415
rect 617 18381 814 18386
rect 848 18381 1026 18415
rect 617 18352 1026 18381
rect 617 18318 646 18352
rect 680 18343 1026 18352
rect 680 18318 814 18343
rect 617 18309 814 18318
rect 848 18309 1026 18343
rect 617 18284 1026 18309
rect 617 18250 646 18284
rect 680 18271 1026 18284
rect 680 18250 814 18271
rect 617 18237 814 18250
rect 848 18237 1026 18271
rect 617 18216 1026 18237
rect 617 18182 646 18216
rect 680 18199 1026 18216
rect 680 18182 814 18199
rect 617 18165 814 18182
rect 848 18165 1026 18199
rect 617 18148 1026 18165
rect 617 18114 646 18148
rect 680 18127 1026 18148
rect 680 18114 814 18127
rect 617 18093 814 18114
rect 848 18093 1026 18127
rect 617 18080 1026 18093
rect 617 18046 646 18080
rect 680 18055 1026 18080
rect 680 18046 814 18055
rect 617 18021 814 18046
rect 848 18021 1026 18055
rect 617 18012 1026 18021
rect 617 17978 646 18012
rect 680 17983 1026 18012
rect 680 17978 814 17983
rect 617 17949 814 17978
rect 848 17949 1026 17983
rect 617 17944 1026 17949
rect 617 17910 646 17944
rect 680 17911 1026 17944
rect 680 17910 814 17911
rect 617 17877 814 17910
rect 848 17877 1026 17911
rect 617 17876 1026 17877
rect 617 17842 646 17876
rect 680 17842 1026 17876
rect 617 17839 1026 17842
rect 617 17808 814 17839
rect 617 17774 646 17808
rect 680 17805 814 17808
rect 848 17805 1026 17839
rect 680 17774 1026 17805
rect 617 17767 1026 17774
rect 617 17740 814 17767
rect 617 17706 646 17740
rect 680 17733 814 17740
rect 848 17733 1026 17767
rect 680 17706 1026 17733
rect 617 17695 1026 17706
rect 617 17672 814 17695
rect 617 17638 646 17672
rect 680 17661 814 17672
rect 848 17661 1026 17695
rect 680 17638 1026 17661
rect 617 17623 1026 17638
rect 617 17604 814 17623
rect 617 17570 646 17604
rect 680 17589 814 17604
rect 848 17589 1026 17623
rect 680 17570 1026 17589
rect 617 17551 1026 17570
rect 617 17536 814 17551
rect 617 17502 646 17536
rect 680 17517 814 17536
rect 848 17517 1026 17551
rect 680 17502 1026 17517
rect 617 17479 1026 17502
rect 617 17468 814 17479
rect 617 17434 646 17468
rect 680 17445 814 17468
rect 848 17445 1026 17479
rect 680 17434 1026 17445
rect 617 17407 1026 17434
rect 617 17400 814 17407
rect 617 17366 646 17400
rect 680 17373 814 17400
rect 848 17373 1026 17407
rect 680 17366 1026 17373
rect 617 17335 1026 17366
rect 617 17332 814 17335
rect 617 17298 646 17332
rect 680 17301 814 17332
rect 848 17301 1026 17335
rect 680 17298 1026 17301
rect 617 17264 1026 17298
rect 617 17230 646 17264
rect 680 17263 1026 17264
rect 680 17230 814 17263
rect 617 17229 814 17230
rect 848 17229 1026 17263
rect 617 17196 1026 17229
rect 617 17162 646 17196
rect 680 17191 1026 17196
rect 680 17162 814 17191
rect 617 17157 814 17162
rect 848 17157 1026 17191
rect 617 17128 1026 17157
rect 617 17094 646 17128
rect 680 17119 1026 17128
rect 680 17094 814 17119
rect 617 17085 814 17094
rect 848 17085 1026 17119
rect 617 17060 1026 17085
rect 617 17026 646 17060
rect 680 17047 1026 17060
rect 680 17026 814 17047
rect 617 17013 814 17026
rect 848 17013 1026 17047
rect 617 16992 1026 17013
rect 617 16958 646 16992
rect 680 16975 1026 16992
rect 680 16958 814 16975
rect 617 16941 814 16958
rect 848 16941 1026 16975
rect 617 16924 1026 16941
rect 617 16890 646 16924
rect 680 16903 1026 16924
rect 680 16890 814 16903
rect 617 16869 814 16890
rect 848 16869 1026 16903
rect 617 16856 1026 16869
rect 617 16822 646 16856
rect 680 16831 1026 16856
rect 680 16822 814 16831
rect 617 16797 814 16822
rect 848 16797 1026 16831
rect 617 16788 1026 16797
rect 617 16754 646 16788
rect 680 16759 1026 16788
rect 680 16754 814 16759
rect 617 16725 814 16754
rect 848 16725 1026 16759
rect 617 16720 1026 16725
rect 617 16686 646 16720
rect 680 16687 1026 16720
rect 680 16686 814 16687
rect 617 16653 814 16686
rect 848 16653 1026 16687
rect 617 16652 1026 16653
rect 617 16618 646 16652
rect 680 16618 1026 16652
rect 617 16615 1026 16618
rect 617 16584 814 16615
rect 617 16550 646 16584
rect 680 16581 814 16584
rect 848 16581 1026 16615
rect 680 16550 1026 16581
rect 617 16543 1026 16550
rect 617 16516 814 16543
rect 617 16482 646 16516
rect 680 16509 814 16516
rect 848 16509 1026 16543
rect 680 16482 1026 16509
rect 617 16471 1026 16482
rect 617 16448 814 16471
rect 617 16414 646 16448
rect 680 16437 814 16448
rect 848 16437 1026 16471
rect 680 16414 1026 16437
rect 617 16399 1026 16414
rect 617 16380 814 16399
rect 617 16346 646 16380
rect 680 16365 814 16380
rect 848 16365 1026 16399
rect 680 16346 1026 16365
rect 617 16327 1026 16346
rect 617 16312 814 16327
rect 617 16278 646 16312
rect 680 16293 814 16312
rect 848 16293 1026 16327
rect 680 16278 1026 16293
rect 617 16255 1026 16278
rect 617 16244 814 16255
rect 617 16210 646 16244
rect 680 16221 814 16244
rect 848 16221 1026 16255
rect 680 16210 1026 16221
rect 617 16183 1026 16210
rect 617 16176 814 16183
rect 617 16142 646 16176
rect 680 16149 814 16176
rect 848 16149 1026 16183
rect 680 16142 1026 16149
rect 617 16111 1026 16142
rect 617 16108 814 16111
rect 617 16074 646 16108
rect 680 16077 814 16108
rect 848 16077 1026 16111
rect 680 16074 1026 16077
rect 617 16040 1026 16074
rect 617 16006 646 16040
rect 680 16039 1026 16040
rect 680 16006 814 16039
rect 617 16005 814 16006
rect 848 16005 1026 16039
rect 617 15972 1026 16005
rect 617 15938 646 15972
rect 680 15967 1026 15972
rect 680 15938 814 15967
rect 617 15933 814 15938
rect 848 15933 1026 15967
rect 617 15904 1026 15933
rect 617 15870 646 15904
rect 680 15895 1026 15904
rect 680 15870 814 15895
rect 617 15861 814 15870
rect 848 15861 1026 15895
rect 617 15836 1026 15861
rect 617 15802 646 15836
rect 680 15823 1026 15836
rect 680 15802 814 15823
rect 617 15789 814 15802
rect 848 15789 1026 15823
rect 617 15768 1026 15789
rect 617 15734 646 15768
rect 680 15751 1026 15768
rect 680 15734 814 15751
rect 617 15717 814 15734
rect 848 15717 1026 15751
rect 617 15700 1026 15717
rect 617 15666 646 15700
rect 680 15679 1026 15700
rect 680 15666 814 15679
rect 617 15645 814 15666
rect 848 15645 1026 15679
rect 617 15632 1026 15645
rect 617 15598 646 15632
rect 680 15607 1026 15632
rect 680 15598 814 15607
rect 617 15573 814 15598
rect 848 15573 1026 15607
rect 617 15564 1026 15573
rect 617 15530 646 15564
rect 680 15535 1026 15564
rect 680 15530 814 15535
rect 617 15501 814 15530
rect 848 15501 1026 15535
rect 617 15496 1026 15501
rect 617 15462 646 15496
rect 680 15463 1026 15496
rect 680 15462 814 15463
rect 617 15429 814 15462
rect 848 15429 1026 15463
rect 617 15428 1026 15429
rect 617 15394 646 15428
rect 680 15394 1026 15428
rect 617 15391 1026 15394
rect 617 15360 814 15391
rect 617 15326 646 15360
rect 680 15357 814 15360
rect 848 15357 1026 15391
rect 680 15326 1026 15357
rect 617 15319 1026 15326
rect 617 15292 814 15319
rect 617 15258 646 15292
rect 680 15285 814 15292
rect 848 15285 1026 15319
rect 680 15258 1026 15285
rect 617 15247 1026 15258
rect 617 15224 814 15247
rect 617 15190 646 15224
rect 680 15213 814 15224
rect 848 15213 1026 15247
rect 680 15190 1026 15213
rect 617 15175 1026 15190
rect 617 15156 814 15175
rect 617 15122 646 15156
rect 680 15141 814 15156
rect 848 15141 1026 15175
rect 680 15122 1026 15141
rect 617 15103 1026 15122
rect 617 15088 814 15103
rect 617 15054 646 15088
rect 680 15069 814 15088
rect 848 15069 1026 15103
rect 680 15054 1026 15069
rect 617 15031 1026 15054
rect 617 15020 814 15031
rect 617 14986 646 15020
rect 680 14997 814 15020
rect 848 14997 1026 15031
rect 680 14986 1026 14997
rect 617 14959 1026 14986
rect 617 14952 814 14959
rect 617 14918 646 14952
rect 680 14925 814 14952
rect 848 14925 1026 14959
rect 680 14918 1026 14925
rect 617 14887 1026 14918
rect 617 14884 814 14887
rect 617 14850 646 14884
rect 680 14853 814 14884
rect 848 14853 1026 14887
rect 680 14850 1026 14853
rect 617 14816 1026 14850
rect 617 14782 646 14816
rect 680 14815 1026 14816
rect 680 14782 814 14815
rect 617 14781 814 14782
rect 848 14781 1026 14815
rect 617 14748 1026 14781
rect 617 14714 646 14748
rect 680 14743 1026 14748
rect 680 14714 814 14743
rect 617 14709 814 14714
rect 848 14709 1026 14743
rect 617 14680 1026 14709
rect 617 14646 646 14680
rect 680 14671 1026 14680
rect 680 14646 814 14671
rect 617 14637 814 14646
rect 848 14637 1026 14671
rect 617 14612 1026 14637
rect 617 14578 646 14612
rect 680 14599 1026 14612
rect 680 14578 814 14599
rect 617 14565 814 14578
rect 848 14565 1026 14599
rect 617 14544 1026 14565
rect 617 14510 646 14544
rect 680 14527 1026 14544
rect 680 14510 814 14527
rect 617 14493 814 14510
rect 848 14493 1026 14527
rect 617 14476 1026 14493
rect 617 14442 646 14476
rect 680 14455 1026 14476
rect 680 14442 814 14455
rect 617 14421 814 14442
rect 848 14421 1026 14455
rect 617 14408 1026 14421
rect 617 14374 646 14408
rect 680 14383 1026 14408
rect 680 14374 814 14383
rect 617 14349 814 14374
rect 848 14349 1026 14383
rect 617 14340 1026 14349
rect 617 14306 646 14340
rect 680 14311 1026 14340
rect 680 14306 814 14311
rect 617 14277 814 14306
rect 848 14277 1026 14311
rect 617 14272 1026 14277
rect 617 14238 646 14272
rect 680 14239 1026 14272
rect 680 14238 814 14239
rect 617 14205 814 14238
rect 848 14205 1026 14239
rect 617 14204 1026 14205
rect 617 14170 646 14204
rect 680 14170 1026 14204
rect 617 14167 1026 14170
rect 617 14136 814 14167
rect 617 14102 646 14136
rect 680 14133 814 14136
rect 848 14133 1026 14167
rect 680 14102 1026 14133
rect 617 14095 1026 14102
rect 617 14068 814 14095
rect 617 14034 646 14068
rect 680 14061 814 14068
rect 848 14061 1026 14095
rect 680 14034 1026 14061
rect 617 14023 1026 14034
rect 617 14000 814 14023
rect 617 13966 646 14000
rect 680 13989 814 14000
rect 848 13989 1026 14023
rect 680 13966 1026 13989
rect 617 13951 1026 13966
rect 617 13932 814 13951
rect 617 13898 646 13932
rect 680 13917 814 13932
rect 848 13917 1026 13951
rect 680 13898 1026 13917
rect 617 13879 1026 13898
rect 617 13864 814 13879
rect 617 13830 646 13864
rect 680 13845 814 13864
rect 848 13845 1026 13879
rect 680 13830 1026 13845
rect 617 13807 1026 13830
rect 617 13796 814 13807
rect 617 13762 646 13796
rect 680 13773 814 13796
rect 848 13773 1026 13807
rect 680 13762 1026 13773
rect 617 13735 1026 13762
rect 617 13728 814 13735
rect 617 13694 646 13728
rect 680 13701 814 13728
rect 848 13701 1026 13735
rect 680 13694 1026 13701
rect 617 13663 1026 13694
rect 617 13660 814 13663
rect 617 13626 646 13660
rect 680 13629 814 13660
rect 848 13629 1026 13663
rect 680 13626 1026 13629
rect 617 13592 1026 13626
rect 617 13558 646 13592
rect 680 13591 1026 13592
rect 680 13558 814 13591
rect 617 13557 814 13558
rect 848 13557 1026 13591
rect 617 13524 1026 13557
rect 617 13490 646 13524
rect 680 13519 1026 13524
rect 680 13490 814 13519
rect 617 13485 814 13490
rect 848 13485 1026 13519
rect 617 13456 1026 13485
rect 617 13422 646 13456
rect 680 13447 1026 13456
rect 680 13422 814 13447
rect 617 13413 814 13422
rect 848 13413 1026 13447
rect 617 13388 1026 13413
rect 617 13354 646 13388
rect 680 13375 1026 13388
rect 680 13354 814 13375
rect 617 13341 814 13354
rect 848 13341 1026 13375
rect 617 13320 1026 13341
rect 617 13286 646 13320
rect 680 13303 1026 13320
rect 680 13286 814 13303
rect 617 13269 814 13286
rect 848 13269 1026 13303
rect 617 13252 1026 13269
rect 617 13218 646 13252
rect 680 13231 1026 13252
rect 680 13218 814 13231
rect 617 13197 814 13218
rect 848 13197 1026 13231
rect 617 13184 1026 13197
rect 617 13150 646 13184
rect 680 13159 1026 13184
rect 680 13150 814 13159
rect 617 13125 814 13150
rect 848 13125 1026 13159
rect 617 13116 1026 13125
rect 617 13082 646 13116
rect 680 13087 1026 13116
rect 680 13082 814 13087
rect 617 13053 814 13082
rect 848 13053 1026 13087
rect 617 13048 1026 13053
rect 617 13014 646 13048
rect 680 13015 1026 13048
rect 680 13014 814 13015
rect 617 12981 814 13014
rect 848 12981 1026 13015
rect 617 12980 1026 12981
rect 617 12946 646 12980
rect 680 12946 1026 12980
rect 617 12943 1026 12946
rect 617 12912 814 12943
rect 617 12878 646 12912
rect 680 12909 814 12912
rect 848 12909 1026 12943
rect 680 12878 1026 12909
rect 617 12871 1026 12878
rect 617 12844 814 12871
rect 617 12810 646 12844
rect 680 12837 814 12844
rect 848 12837 1026 12871
rect 680 12810 1026 12837
rect 617 12799 1026 12810
rect 617 12776 814 12799
rect 617 12742 646 12776
rect 680 12765 814 12776
rect 848 12765 1026 12799
rect 680 12742 1026 12765
rect 617 12727 1026 12742
rect 617 12708 814 12727
rect 617 12674 646 12708
rect 680 12693 814 12708
rect 848 12693 1026 12727
rect 680 12674 1026 12693
rect 617 12655 1026 12674
rect 617 12640 814 12655
rect 617 12606 646 12640
rect 680 12621 814 12640
rect 848 12621 1026 12655
rect 680 12606 1026 12621
rect 617 12583 1026 12606
rect 617 12572 814 12583
rect 617 12538 646 12572
rect 680 12549 814 12572
rect 848 12549 1026 12583
rect 680 12538 1026 12549
rect 617 12511 1026 12538
rect 617 12504 814 12511
rect 617 12470 646 12504
rect 680 12477 814 12504
rect 848 12477 1026 12511
rect 680 12470 1026 12477
rect 617 12439 1026 12470
rect 617 12436 814 12439
rect 617 12402 646 12436
rect 680 12405 814 12436
rect 848 12405 1026 12439
rect 680 12402 1026 12405
rect 617 12368 1026 12402
rect 617 12334 646 12368
rect 680 12367 1026 12368
rect 680 12334 814 12367
rect 617 12333 814 12334
rect 848 12333 1026 12367
rect 617 12300 1026 12333
rect 617 12266 646 12300
rect 680 12295 1026 12300
rect 680 12266 814 12295
rect 617 12261 814 12266
rect 848 12261 1026 12295
rect 617 12232 1026 12261
rect 617 12198 646 12232
rect 680 12223 1026 12232
rect 680 12198 814 12223
rect 617 12189 814 12198
rect 848 12189 1026 12223
rect 617 12164 1026 12189
rect 617 12130 646 12164
rect 680 12151 1026 12164
rect 680 12130 814 12151
rect 617 12117 814 12130
rect 848 12117 1026 12151
rect 617 12096 1026 12117
rect 617 12062 646 12096
rect 680 12079 1026 12096
rect 680 12062 814 12079
rect 617 12045 814 12062
rect 848 12045 1026 12079
rect 617 12028 1026 12045
rect 617 11994 646 12028
rect 680 12007 1026 12028
rect 680 11994 814 12007
rect 617 11973 814 11994
rect 848 11973 1026 12007
rect 617 11960 1026 11973
rect 617 11926 646 11960
rect 680 11935 1026 11960
rect 680 11926 814 11935
rect 617 11901 814 11926
rect 848 11901 1026 11935
rect 617 11892 1026 11901
rect 617 11858 646 11892
rect 680 11863 1026 11892
rect 680 11858 814 11863
rect 617 11829 814 11858
rect 848 11829 1026 11863
rect 617 11824 1026 11829
rect 617 11790 646 11824
rect 680 11791 1026 11824
rect 680 11790 814 11791
rect 617 11757 814 11790
rect 848 11757 1026 11791
rect 617 11756 1026 11757
rect 617 11722 646 11756
rect 680 11722 1026 11756
rect 617 11719 1026 11722
rect 617 11688 814 11719
rect 617 11654 646 11688
rect 680 11685 814 11688
rect 848 11685 1026 11719
rect 680 11654 1026 11685
rect 617 11647 1026 11654
rect 617 11620 814 11647
rect 617 11586 646 11620
rect 680 11613 814 11620
rect 848 11613 1026 11647
rect 680 11586 1026 11613
rect 617 11575 1026 11586
rect 617 11552 814 11575
rect 617 11518 646 11552
rect 680 11541 814 11552
rect 848 11541 1026 11575
rect 680 11518 1026 11541
rect 617 11503 1026 11518
rect 617 11484 814 11503
rect 617 11450 646 11484
rect 680 11469 814 11484
rect 848 11469 1026 11503
rect 680 11450 1026 11469
rect 617 11431 1026 11450
rect 617 11416 814 11431
rect 617 11382 646 11416
rect 680 11397 814 11416
rect 848 11397 1026 11431
rect 680 11382 1026 11397
rect 617 11359 1026 11382
rect 617 11348 814 11359
rect 617 11314 646 11348
rect 680 11325 814 11348
rect 848 11325 1026 11359
rect 680 11314 1026 11325
rect 617 11287 1026 11314
rect 617 11280 814 11287
rect 617 11246 646 11280
rect 680 11253 814 11280
rect 848 11253 1026 11287
rect 680 11246 1026 11253
rect 617 11215 1026 11246
rect 617 11212 814 11215
rect 617 11178 646 11212
rect 680 11181 814 11212
rect 848 11181 1026 11215
rect 680 11178 1026 11181
rect 617 11144 1026 11178
rect 617 11110 646 11144
rect 680 11143 1026 11144
rect 680 11110 814 11143
rect 617 11109 814 11110
rect 848 11109 1026 11143
rect 617 11076 1026 11109
rect 617 11042 646 11076
rect 680 11071 1026 11076
rect 680 11042 814 11071
rect 617 11037 814 11042
rect 848 11037 1026 11071
rect 617 11008 1026 11037
rect 617 10974 646 11008
rect 680 10999 1026 11008
rect 680 10974 814 10999
rect 617 10965 814 10974
rect 848 10965 1026 10999
rect 617 10940 1026 10965
rect 617 10906 646 10940
rect 680 10927 1026 10940
rect 680 10906 814 10927
rect 617 10893 814 10906
rect 848 10893 1026 10927
rect 617 10872 1026 10893
rect 617 10838 646 10872
rect 680 10855 1026 10872
rect 680 10838 814 10855
rect 617 10821 814 10838
rect 848 10821 1026 10855
rect 617 10804 1026 10821
rect 617 10770 646 10804
rect 680 10783 1026 10804
rect 680 10770 814 10783
rect 617 10749 814 10770
rect 848 10749 1026 10783
rect 617 10736 1026 10749
rect 617 10702 646 10736
rect 680 10711 1026 10736
rect 680 10702 814 10711
rect 617 10677 814 10702
rect 848 10677 1026 10711
rect 617 10668 1026 10677
rect 617 10634 646 10668
rect 680 10639 1026 10668
rect 680 10634 814 10639
rect 617 10605 814 10634
rect 848 10605 1026 10639
rect 617 10600 1026 10605
rect 617 10566 646 10600
rect 680 10567 1026 10600
rect 680 10566 814 10567
rect 617 10533 814 10566
rect 848 10533 1026 10567
rect 617 10532 1026 10533
rect 617 10498 646 10532
rect 680 10498 1026 10532
rect 617 10495 1026 10498
rect 617 10464 814 10495
rect 617 10430 646 10464
rect 680 10461 814 10464
rect 848 10461 1026 10495
rect 680 10430 1026 10461
rect 617 10423 1026 10430
rect 617 10396 814 10423
rect 617 10362 646 10396
rect 680 10389 814 10396
rect 848 10389 1026 10423
rect 680 10362 1026 10389
rect 617 10351 1026 10362
rect 617 10328 814 10351
rect 617 10294 646 10328
rect 680 10317 814 10328
rect 848 10317 1026 10351
rect 680 10294 1026 10317
rect 617 10279 1026 10294
rect 617 10260 814 10279
rect 617 10226 646 10260
rect 680 10245 814 10260
rect 848 10245 1026 10279
rect 680 10226 1026 10245
rect 617 10207 1026 10226
rect 1177 34636 13817 34684
rect 1177 34602 1365 34636
rect 1399 34602 1433 34636
rect 1471 34602 1501 34636
rect 1543 34602 1569 34636
rect 1615 34602 1637 34636
rect 1687 34602 1705 34636
rect 1759 34602 1773 34636
rect 1831 34602 1841 34636
rect 1903 34602 1909 34636
rect 1975 34602 1977 34636
rect 2011 34602 2013 34636
rect 2079 34602 2085 34636
rect 2147 34602 2157 34636
rect 2215 34602 2229 34636
rect 2283 34602 2301 34636
rect 2351 34602 2373 34636
rect 2419 34602 2445 34636
rect 2487 34602 2517 34636
rect 2555 34602 2589 34636
rect 2623 34602 2657 34636
rect 2695 34602 2725 34636
rect 2767 34602 2793 34636
rect 2839 34602 2861 34636
rect 2911 34602 2929 34636
rect 2983 34602 2997 34636
rect 3055 34602 3065 34636
rect 3127 34602 3133 34636
rect 3199 34602 3201 34636
rect 3235 34602 3237 34636
rect 3303 34602 3309 34636
rect 3371 34602 3381 34636
rect 3439 34602 3453 34636
rect 3507 34602 3525 34636
rect 3575 34602 3597 34636
rect 3643 34602 3669 34636
rect 3711 34602 3741 34636
rect 3779 34602 3813 34636
rect 3847 34602 3881 34636
rect 3919 34602 3949 34636
rect 3991 34602 4017 34636
rect 4063 34602 4085 34636
rect 4135 34602 4153 34636
rect 4207 34602 4221 34636
rect 4279 34602 4289 34636
rect 4351 34602 4357 34636
rect 4423 34602 4425 34636
rect 4459 34602 4461 34636
rect 4527 34602 4533 34636
rect 4595 34602 4605 34636
rect 4663 34602 4677 34636
rect 4731 34602 4749 34636
rect 4799 34602 4821 34636
rect 4867 34602 4893 34636
rect 4935 34602 4965 34636
rect 5003 34602 5037 34636
rect 5071 34602 5105 34636
rect 5143 34602 5173 34636
rect 5215 34602 5241 34636
rect 5287 34602 5309 34636
rect 5359 34602 5377 34636
rect 5431 34602 5445 34636
rect 5503 34602 5513 34636
rect 5575 34602 5581 34636
rect 5647 34602 5649 34636
rect 5683 34602 5685 34636
rect 5751 34602 5757 34636
rect 5819 34602 5829 34636
rect 5887 34602 5901 34636
rect 5955 34602 5973 34636
rect 6023 34602 6045 34636
rect 6091 34602 6117 34636
rect 6159 34602 6189 34636
rect 6227 34602 6261 34636
rect 6295 34602 6329 34636
rect 6367 34602 6397 34636
rect 6439 34602 6465 34636
rect 6511 34602 6533 34636
rect 6583 34602 6601 34636
rect 6655 34602 6669 34636
rect 6727 34602 6737 34636
rect 6799 34602 6805 34636
rect 6871 34602 6873 34636
rect 6907 34602 6909 34636
rect 6975 34602 6981 34636
rect 7043 34602 7053 34636
rect 7111 34602 7125 34636
rect 7179 34602 7197 34636
rect 7247 34602 7269 34636
rect 7315 34602 7341 34636
rect 7383 34602 7413 34636
rect 7451 34602 7485 34636
rect 7519 34602 7553 34636
rect 7591 34602 7621 34636
rect 7663 34602 7689 34636
rect 7735 34602 7757 34636
rect 7807 34602 7825 34636
rect 7879 34602 7893 34636
rect 7951 34602 7961 34636
rect 8023 34602 8029 34636
rect 8095 34602 8097 34636
rect 8131 34602 8133 34636
rect 8199 34602 8205 34636
rect 8267 34602 8277 34636
rect 8335 34602 8349 34636
rect 8403 34602 8421 34636
rect 8471 34602 8493 34636
rect 8539 34602 8565 34636
rect 8607 34602 8637 34636
rect 8675 34602 8709 34636
rect 8743 34602 8777 34636
rect 8815 34602 8845 34636
rect 8887 34602 8913 34636
rect 8959 34602 8981 34636
rect 9031 34602 9049 34636
rect 9103 34602 9117 34636
rect 9175 34602 9185 34636
rect 9247 34602 9253 34636
rect 9319 34602 9321 34636
rect 9355 34602 9357 34636
rect 9423 34602 9429 34636
rect 9491 34602 9501 34636
rect 9559 34602 9573 34636
rect 9627 34602 9645 34636
rect 9695 34602 9717 34636
rect 9763 34602 9789 34636
rect 9831 34602 9861 34636
rect 9899 34602 9933 34636
rect 9967 34602 10001 34636
rect 10039 34602 10069 34636
rect 10111 34602 10137 34636
rect 10183 34602 10205 34636
rect 10255 34602 10273 34636
rect 10327 34602 10341 34636
rect 10399 34602 10409 34636
rect 10471 34602 10477 34636
rect 10543 34602 10545 34636
rect 10579 34602 10581 34636
rect 10647 34602 10653 34636
rect 10715 34602 10725 34636
rect 10783 34602 10797 34636
rect 10851 34602 10869 34636
rect 10919 34602 10941 34636
rect 10987 34602 11013 34636
rect 11055 34602 11085 34636
rect 11123 34602 11157 34636
rect 11191 34602 11225 34636
rect 11263 34602 11293 34636
rect 11335 34602 11361 34636
rect 11407 34602 11429 34636
rect 11479 34602 11497 34636
rect 11551 34602 11565 34636
rect 11623 34602 11633 34636
rect 11695 34602 11701 34636
rect 11767 34602 11769 34636
rect 11803 34602 11805 34636
rect 11871 34602 11877 34636
rect 11939 34602 11949 34636
rect 12007 34602 12021 34636
rect 12075 34602 12093 34636
rect 12143 34602 12165 34636
rect 12211 34602 12237 34636
rect 12279 34602 12309 34636
rect 12347 34602 12381 34636
rect 12415 34602 12449 34636
rect 12487 34602 12517 34636
rect 12559 34602 12585 34636
rect 12631 34602 12653 34636
rect 12703 34602 12721 34636
rect 12775 34602 12789 34636
rect 12847 34602 12857 34636
rect 12919 34602 12925 34636
rect 12991 34602 12993 34636
rect 13027 34602 13029 34636
rect 13095 34602 13101 34636
rect 13163 34602 13173 34636
rect 13231 34602 13245 34636
rect 13299 34602 13317 34636
rect 13367 34602 13389 34636
rect 13435 34602 13461 34636
rect 13503 34602 13533 34636
rect 13571 34602 13605 34636
rect 13639 34602 13817 34636
rect 1177 34564 13817 34602
rect 1177 34486 1297 34564
rect 1177 34440 1221 34486
rect 1255 34440 1297 34486
rect 1177 34418 1297 34440
rect 1177 34368 1221 34418
rect 1255 34368 1297 34418
rect 1177 34350 1297 34368
rect 1177 34296 1221 34350
rect 1255 34296 1297 34350
rect 1177 34282 1297 34296
rect 1177 34224 1221 34282
rect 1255 34224 1297 34282
rect 1177 34214 1297 34224
rect 1177 34152 1221 34214
rect 1255 34152 1297 34214
rect 1177 34146 1297 34152
rect 1177 34080 1221 34146
rect 1255 34080 1297 34146
rect 1177 34078 1297 34080
rect 1177 34044 1221 34078
rect 1255 34044 1297 34078
rect 1177 34042 1297 34044
rect 1177 33976 1221 34042
rect 1255 33976 1297 34042
rect 1177 33970 1297 33976
rect 1177 33908 1221 33970
rect 1255 33908 1297 33970
rect 1177 33898 1297 33908
rect 1177 33840 1221 33898
rect 1255 33840 1297 33898
rect 1177 33826 1297 33840
rect 1177 33772 1221 33826
rect 1255 33772 1297 33826
rect 1177 33754 1297 33772
rect 1177 33704 1221 33754
rect 1255 33704 1297 33754
rect 1177 33682 1297 33704
rect 1177 33636 1221 33682
rect 1255 33636 1297 33682
rect 1177 33610 1297 33636
rect 1177 33568 1221 33610
rect 1255 33568 1297 33610
rect 1177 33538 1297 33568
rect 1177 33500 1221 33538
rect 1255 33500 1297 33538
rect 1177 33466 1297 33500
rect 1177 33432 1221 33466
rect 1255 33432 1297 33466
rect 1177 33398 1297 33432
rect 1177 33360 1221 33398
rect 1255 33360 1297 33398
rect 1177 33330 1297 33360
rect 1177 33288 1221 33330
rect 1255 33288 1297 33330
rect 1177 33262 1297 33288
rect 1177 33216 1221 33262
rect 1255 33216 1297 33262
rect 1177 33194 1297 33216
rect 1177 33144 1221 33194
rect 1255 33144 1297 33194
rect 1177 33126 1297 33144
rect 1177 33072 1221 33126
rect 1255 33072 1297 33126
rect 1177 33058 1297 33072
rect 1177 33000 1221 33058
rect 1255 33000 1297 33058
rect 1177 32990 1297 33000
rect 1177 32928 1221 32990
rect 1255 32928 1297 32990
rect 1177 32922 1297 32928
rect 1177 32856 1221 32922
rect 1255 32856 1297 32922
rect 1177 32854 1297 32856
rect 1177 32820 1221 32854
rect 1255 32820 1297 32854
rect 1177 32818 1297 32820
rect 1177 32752 1221 32818
rect 1255 32752 1297 32818
rect 1177 32746 1297 32752
rect 1177 32684 1221 32746
rect 1255 32684 1297 32746
rect 1177 32674 1297 32684
rect 1177 32616 1221 32674
rect 1255 32616 1297 32674
rect 1177 32602 1297 32616
rect 1177 32548 1221 32602
rect 1255 32548 1297 32602
rect 1177 32530 1297 32548
rect 1177 32480 1221 32530
rect 1255 32480 1297 32530
rect 1177 32458 1297 32480
rect 1177 32412 1221 32458
rect 1255 32412 1297 32458
rect 1177 32386 1297 32412
rect 1177 32344 1221 32386
rect 1255 32344 1297 32386
rect 1177 32314 1297 32344
rect 1177 32276 1221 32314
rect 1255 32276 1297 32314
rect 1177 32242 1297 32276
rect 1177 32208 1221 32242
rect 1255 32208 1297 32242
rect 1177 32174 1297 32208
rect 1177 32136 1221 32174
rect 1255 32136 1297 32174
rect 1177 32106 1297 32136
rect 1177 32064 1221 32106
rect 1255 32064 1297 32106
rect 1177 32038 1297 32064
rect 1177 31992 1221 32038
rect 1255 31992 1297 32038
rect 1177 31970 1297 31992
rect 1177 31920 1221 31970
rect 1255 31920 1297 31970
rect 1177 31902 1297 31920
rect 1177 31848 1221 31902
rect 1255 31848 1297 31902
rect 1177 31834 1297 31848
rect 1177 31776 1221 31834
rect 1255 31776 1297 31834
rect 1177 31766 1297 31776
rect 1177 31704 1221 31766
rect 1255 31704 1297 31766
rect 1177 31698 1297 31704
rect 1177 31632 1221 31698
rect 1255 31632 1297 31698
rect 1177 31630 1297 31632
rect 1177 31596 1221 31630
rect 1255 31596 1297 31630
rect 1177 31594 1297 31596
rect 1177 31528 1221 31594
rect 1255 31528 1297 31594
rect 1177 31522 1297 31528
rect 1177 31460 1221 31522
rect 1255 31460 1297 31522
rect 1177 31450 1297 31460
rect 1177 31392 1221 31450
rect 1255 31392 1297 31450
rect 1177 31378 1297 31392
rect 1177 31324 1221 31378
rect 1255 31324 1297 31378
rect 1177 31306 1297 31324
rect 1177 31256 1221 31306
rect 1255 31256 1297 31306
rect 1177 31234 1297 31256
rect 1177 31188 1221 31234
rect 1255 31188 1297 31234
rect 1177 31162 1297 31188
rect 1177 31120 1221 31162
rect 1255 31120 1297 31162
rect 1177 31090 1297 31120
rect 1177 31052 1221 31090
rect 1255 31052 1297 31090
rect 1177 31018 1297 31052
rect 1177 30984 1221 31018
rect 1255 30984 1297 31018
rect 1177 30950 1297 30984
rect 1177 30912 1221 30950
rect 1255 30912 1297 30950
rect 1177 30882 1297 30912
rect 1177 30840 1221 30882
rect 1255 30840 1297 30882
rect 1177 30814 1297 30840
rect 1177 30768 1221 30814
rect 1255 30768 1297 30814
rect 1177 30746 1297 30768
rect 1177 30696 1221 30746
rect 1255 30696 1297 30746
rect 1177 30678 1297 30696
rect 1177 30624 1221 30678
rect 1255 30624 1297 30678
rect 1177 30610 1297 30624
rect 1177 30552 1221 30610
rect 1255 30552 1297 30610
rect 1177 30542 1297 30552
rect 1177 30480 1221 30542
rect 1255 30480 1297 30542
rect 1177 30474 1297 30480
rect 1177 30408 1221 30474
rect 1255 30408 1297 30474
rect 1177 30406 1297 30408
rect 1177 30372 1221 30406
rect 1255 30372 1297 30406
rect 1177 30370 1297 30372
rect 1177 30304 1221 30370
rect 1255 30304 1297 30370
rect 1177 30298 1297 30304
rect 1177 30236 1221 30298
rect 1255 30236 1297 30298
rect 1177 30226 1297 30236
rect 1177 30168 1221 30226
rect 1255 30168 1297 30226
rect 1177 30154 1297 30168
rect 1177 30100 1221 30154
rect 1255 30100 1297 30154
rect 1177 30082 1297 30100
rect 1177 30032 1221 30082
rect 1255 30032 1297 30082
rect 1177 30010 1297 30032
rect 1177 29964 1221 30010
rect 1255 29964 1297 30010
rect 1177 29938 1297 29964
rect 1177 29896 1221 29938
rect 1255 29896 1297 29938
rect 1177 29866 1297 29896
rect 1177 29828 1221 29866
rect 1255 29828 1297 29866
rect 1177 29794 1297 29828
rect 1177 29760 1221 29794
rect 1255 29760 1297 29794
rect 1177 29726 1297 29760
rect 1177 29688 1221 29726
rect 1255 29688 1297 29726
rect 1177 29658 1297 29688
rect 1177 29616 1221 29658
rect 1255 29616 1297 29658
rect 1177 29590 1297 29616
rect 1177 29544 1221 29590
rect 1255 29544 1297 29590
rect 1177 29522 1297 29544
rect 1177 29472 1221 29522
rect 1255 29472 1297 29522
rect 1177 29454 1297 29472
rect 1177 29400 1221 29454
rect 1255 29400 1297 29454
rect 1177 29386 1297 29400
rect 1177 29328 1221 29386
rect 1255 29328 1297 29386
rect 1177 29318 1297 29328
rect 1177 29256 1221 29318
rect 1255 29256 1297 29318
rect 1177 29250 1297 29256
rect 1177 29184 1221 29250
rect 1255 29184 1297 29250
rect 1177 29182 1297 29184
rect 1177 29148 1221 29182
rect 1255 29148 1297 29182
rect 1177 29146 1297 29148
rect 1177 29080 1221 29146
rect 1255 29080 1297 29146
rect 1177 29074 1297 29080
rect 1177 29012 1221 29074
rect 1255 29012 1297 29074
rect 1177 29002 1297 29012
rect 1177 28944 1221 29002
rect 1255 28944 1297 29002
rect 1177 28930 1297 28944
rect 1177 28876 1221 28930
rect 1255 28876 1297 28930
rect 1177 28858 1297 28876
rect 1177 28808 1221 28858
rect 1255 28808 1297 28858
rect 1177 28786 1297 28808
rect 1177 28740 1221 28786
rect 1255 28740 1297 28786
rect 1177 28714 1297 28740
rect 1177 28672 1221 28714
rect 1255 28672 1297 28714
rect 1177 28642 1297 28672
rect 1177 28604 1221 28642
rect 1255 28604 1297 28642
rect 1177 28570 1297 28604
rect 1177 28536 1221 28570
rect 1255 28536 1297 28570
rect 1177 28502 1297 28536
rect 1177 28464 1221 28502
rect 1255 28464 1297 28502
rect 1177 28434 1297 28464
rect 1177 28392 1221 28434
rect 1255 28392 1297 28434
rect 1177 28366 1297 28392
rect 1177 28320 1221 28366
rect 1255 28320 1297 28366
rect 1177 28298 1297 28320
rect 1177 28248 1221 28298
rect 1255 28248 1297 28298
rect 1177 28230 1297 28248
rect 1177 28176 1221 28230
rect 1255 28176 1297 28230
rect 1177 28162 1297 28176
rect 1177 28104 1221 28162
rect 1255 28104 1297 28162
rect 1177 28094 1297 28104
rect 1177 28032 1221 28094
rect 1255 28032 1297 28094
rect 1177 28026 1297 28032
rect 1177 27960 1221 28026
rect 1255 27960 1297 28026
rect 1177 27958 1297 27960
rect 1177 27924 1221 27958
rect 1255 27924 1297 27958
rect 1177 27922 1297 27924
rect 1177 27856 1221 27922
rect 1255 27856 1297 27922
rect 1177 27850 1297 27856
rect 1177 27788 1221 27850
rect 1255 27788 1297 27850
rect 1177 27778 1297 27788
rect 1177 27720 1221 27778
rect 1255 27720 1297 27778
rect 1177 27706 1297 27720
rect 1177 27652 1221 27706
rect 1255 27652 1297 27706
rect 1177 27634 1297 27652
rect 1177 27584 1221 27634
rect 1255 27584 1297 27634
rect 1177 27562 1297 27584
rect 1177 27516 1221 27562
rect 1255 27516 1297 27562
rect 1177 27490 1297 27516
rect 1177 27448 1221 27490
rect 1255 27448 1297 27490
rect 1177 27418 1297 27448
rect 1177 27380 1221 27418
rect 1255 27380 1297 27418
rect 1177 27346 1297 27380
rect 1177 27312 1221 27346
rect 1255 27312 1297 27346
rect 1177 27278 1297 27312
rect 1177 27240 1221 27278
rect 1255 27240 1297 27278
rect 1177 27210 1297 27240
rect 1177 27168 1221 27210
rect 1255 27168 1297 27210
rect 1177 27142 1297 27168
rect 1177 27096 1221 27142
rect 1255 27096 1297 27142
rect 1177 27074 1297 27096
rect 1177 27024 1221 27074
rect 1255 27024 1297 27074
rect 1177 27006 1297 27024
rect 1177 26952 1221 27006
rect 1255 26952 1297 27006
rect 1177 26938 1297 26952
rect 1177 26880 1221 26938
rect 1255 26880 1297 26938
rect 1177 26870 1297 26880
rect 1177 26808 1221 26870
rect 1255 26808 1297 26870
rect 1177 26802 1297 26808
rect 1177 26736 1221 26802
rect 1255 26736 1297 26802
rect 1177 26734 1297 26736
rect 1177 26700 1221 26734
rect 1255 26700 1297 26734
rect 1177 26698 1297 26700
rect 1177 26632 1221 26698
rect 1255 26632 1297 26698
rect 1177 26626 1297 26632
rect 1177 26564 1221 26626
rect 1255 26564 1297 26626
rect 1177 26554 1297 26564
rect 1177 26496 1221 26554
rect 1255 26496 1297 26554
rect 1177 26482 1297 26496
rect 1177 26428 1221 26482
rect 1255 26428 1297 26482
rect 1177 26410 1297 26428
rect 1177 26360 1221 26410
rect 1255 26360 1297 26410
rect 1177 26338 1297 26360
rect 1177 26292 1221 26338
rect 1255 26292 1297 26338
rect 1177 26266 1297 26292
rect 1177 26224 1221 26266
rect 1255 26224 1297 26266
rect 1177 26194 1297 26224
rect 1177 26156 1221 26194
rect 1255 26156 1297 26194
rect 1177 26122 1297 26156
rect 1177 26088 1221 26122
rect 1255 26088 1297 26122
rect 1177 26054 1297 26088
rect 1177 26016 1221 26054
rect 1255 26016 1297 26054
rect 1177 25986 1297 26016
rect 1177 25944 1221 25986
rect 1255 25944 1297 25986
rect 1177 25918 1297 25944
rect 1177 25872 1221 25918
rect 1255 25872 1297 25918
rect 1177 25850 1297 25872
rect 1177 25800 1221 25850
rect 1255 25800 1297 25850
rect 1177 25782 1297 25800
rect 1177 25728 1221 25782
rect 1255 25728 1297 25782
rect 1177 25714 1297 25728
rect 1177 25656 1221 25714
rect 1255 25656 1297 25714
rect 1177 25646 1297 25656
rect 1177 25584 1221 25646
rect 1255 25584 1297 25646
rect 1177 25578 1297 25584
rect 1177 25512 1221 25578
rect 1255 25512 1297 25578
rect 1177 25510 1297 25512
rect 1177 25476 1221 25510
rect 1255 25476 1297 25510
rect 1177 25474 1297 25476
rect 1177 25408 1221 25474
rect 1255 25408 1297 25474
rect 1177 25402 1297 25408
rect 1177 25340 1221 25402
rect 1255 25340 1297 25402
rect 1177 25330 1297 25340
rect 1177 25272 1221 25330
rect 1255 25272 1297 25330
rect 1177 25258 1297 25272
rect 1177 25204 1221 25258
rect 1255 25204 1297 25258
rect 1177 25186 1297 25204
rect 1177 25136 1221 25186
rect 1255 25136 1297 25186
rect 1177 25114 1297 25136
rect 1177 25068 1221 25114
rect 1255 25068 1297 25114
rect 1177 25042 1297 25068
rect 1177 25000 1221 25042
rect 1255 25000 1297 25042
rect 1177 24970 1297 25000
rect 1177 24932 1221 24970
rect 1255 24932 1297 24970
rect 1177 24898 1297 24932
rect 1177 24864 1221 24898
rect 1255 24864 1297 24898
rect 1177 24830 1297 24864
rect 1177 24792 1221 24830
rect 1255 24792 1297 24830
rect 1177 24762 1297 24792
rect 1177 24720 1221 24762
rect 1255 24720 1297 24762
rect 1177 24694 1297 24720
rect 1177 24648 1221 24694
rect 1255 24648 1297 24694
rect 1177 24626 1297 24648
rect 1177 24576 1221 24626
rect 1255 24576 1297 24626
rect 1177 24558 1297 24576
rect 1177 24504 1221 24558
rect 1255 24504 1297 24558
rect 1177 24490 1297 24504
rect 1177 24432 1221 24490
rect 1255 24432 1297 24490
rect 1177 24422 1297 24432
rect 1177 24360 1221 24422
rect 1255 24360 1297 24422
rect 1177 24354 1297 24360
rect 1177 24288 1221 24354
rect 1255 24288 1297 24354
rect 1177 24286 1297 24288
rect 1177 24252 1221 24286
rect 1255 24252 1297 24286
rect 1177 24250 1297 24252
rect 1177 24184 1221 24250
rect 1255 24184 1297 24250
rect 1177 24178 1297 24184
rect 1177 24116 1221 24178
rect 1255 24116 1297 24178
rect 1177 24106 1297 24116
rect 1177 24048 1221 24106
rect 1255 24048 1297 24106
rect 1177 24034 1297 24048
rect 1177 23980 1221 24034
rect 1255 23980 1297 24034
rect 1177 23962 1297 23980
rect 1177 23912 1221 23962
rect 1255 23912 1297 23962
rect 1177 23890 1297 23912
rect 1177 23844 1221 23890
rect 1255 23844 1297 23890
rect 1177 23818 1297 23844
rect 1177 23776 1221 23818
rect 1255 23776 1297 23818
rect 1177 23746 1297 23776
rect 1177 23708 1221 23746
rect 1255 23708 1297 23746
rect 1177 23674 1297 23708
rect 1177 23640 1221 23674
rect 1255 23640 1297 23674
rect 1177 23606 1297 23640
rect 1177 23568 1221 23606
rect 1255 23568 1297 23606
rect 1177 23538 1297 23568
rect 1177 23496 1221 23538
rect 1255 23496 1297 23538
rect 1177 23470 1297 23496
rect 1177 23424 1221 23470
rect 1255 23424 1297 23470
rect 1177 23402 1297 23424
rect 1177 23352 1221 23402
rect 1255 23352 1297 23402
rect 1177 23334 1297 23352
rect 1177 23280 1221 23334
rect 1255 23280 1297 23334
rect 1177 23266 1297 23280
rect 1177 23208 1221 23266
rect 1255 23208 1297 23266
rect 1177 23198 1297 23208
rect 1177 23136 1221 23198
rect 1255 23136 1297 23198
rect 1177 23130 1297 23136
rect 1177 23064 1221 23130
rect 1255 23064 1297 23130
rect 1177 23062 1297 23064
rect 1177 23028 1221 23062
rect 1255 23028 1297 23062
rect 1177 23026 1297 23028
rect 1177 22960 1221 23026
rect 1255 22960 1297 23026
rect 1177 22954 1297 22960
rect 1177 22892 1221 22954
rect 1255 22892 1297 22954
rect 1177 22882 1297 22892
rect 1177 22824 1221 22882
rect 1255 22824 1297 22882
rect 1177 22810 1297 22824
rect 1177 22756 1221 22810
rect 1255 22756 1297 22810
rect 1177 22738 1297 22756
rect 1177 22688 1221 22738
rect 1255 22688 1297 22738
rect 1177 22666 1297 22688
rect 1177 22620 1221 22666
rect 1255 22620 1297 22666
rect 1177 22594 1297 22620
rect 1177 22552 1221 22594
rect 1255 22552 1297 22594
rect 1177 22522 1297 22552
rect 1177 22484 1221 22522
rect 1255 22484 1297 22522
rect 1177 22450 1297 22484
rect 1177 22416 1221 22450
rect 1255 22416 1297 22450
rect 1177 22382 1297 22416
rect 1177 22344 1221 22382
rect 1255 22344 1297 22382
rect 1177 22314 1297 22344
rect 1177 22272 1221 22314
rect 1255 22272 1297 22314
rect 1177 22246 1297 22272
rect 1177 22200 1221 22246
rect 1255 22200 1297 22246
rect 1177 22178 1297 22200
rect 1177 22128 1221 22178
rect 1255 22128 1297 22178
rect 1177 22110 1297 22128
rect 1177 22056 1221 22110
rect 1255 22056 1297 22110
rect 1177 22042 1297 22056
rect 1177 21984 1221 22042
rect 1255 21984 1297 22042
rect 1177 21974 1297 21984
rect 1177 21912 1221 21974
rect 1255 21912 1297 21974
rect 1177 21906 1297 21912
rect 1177 21840 1221 21906
rect 1255 21840 1297 21906
rect 1177 21838 1297 21840
rect 1177 21804 1221 21838
rect 1255 21804 1297 21838
rect 1177 21802 1297 21804
rect 1177 21736 1221 21802
rect 1255 21736 1297 21802
rect 1177 21730 1297 21736
rect 1177 21668 1221 21730
rect 1255 21668 1297 21730
rect 1177 21658 1297 21668
rect 1177 21600 1221 21658
rect 1255 21600 1297 21658
rect 1177 21586 1297 21600
rect 1177 21532 1221 21586
rect 1255 21532 1297 21586
rect 1177 21514 1297 21532
rect 1177 21464 1221 21514
rect 1255 21464 1297 21514
rect 1177 21442 1297 21464
rect 1177 21396 1221 21442
rect 1255 21396 1297 21442
rect 1177 21370 1297 21396
rect 1177 21328 1221 21370
rect 1255 21328 1297 21370
rect 1177 21298 1297 21328
rect 1177 21260 1221 21298
rect 1255 21260 1297 21298
rect 1177 21226 1297 21260
rect 1177 21192 1221 21226
rect 1255 21192 1297 21226
rect 1177 21158 1297 21192
rect 1177 21120 1221 21158
rect 1255 21120 1297 21158
rect 1177 21090 1297 21120
rect 1177 21048 1221 21090
rect 1255 21048 1297 21090
rect 1177 21022 1297 21048
rect 1177 20976 1221 21022
rect 1255 20976 1297 21022
rect 1177 20954 1297 20976
rect 1177 20904 1221 20954
rect 1255 20904 1297 20954
rect 1177 20886 1297 20904
rect 1177 20832 1221 20886
rect 1255 20832 1297 20886
rect 1177 20818 1297 20832
rect 1177 20760 1221 20818
rect 1255 20760 1297 20818
rect 1177 20750 1297 20760
rect 1177 20688 1221 20750
rect 1255 20688 1297 20750
rect 1177 20682 1297 20688
rect 1177 20616 1221 20682
rect 1255 20616 1297 20682
rect 1177 20614 1297 20616
rect 1177 20580 1221 20614
rect 1255 20580 1297 20614
rect 1177 20578 1297 20580
rect 1177 20512 1221 20578
rect 1255 20512 1297 20578
rect 1177 20506 1297 20512
rect 1177 20444 1221 20506
rect 1255 20444 1297 20506
rect 1177 20434 1297 20444
rect 1177 20376 1221 20434
rect 1255 20376 1297 20434
rect 1177 20362 1297 20376
rect 1177 20308 1221 20362
rect 1255 20308 1297 20362
rect 1177 20290 1297 20308
rect 1177 20240 1221 20290
rect 1255 20240 1297 20290
rect 1177 20218 1297 20240
rect 1177 20172 1221 20218
rect 1255 20172 1297 20218
rect 1177 20146 1297 20172
rect 1177 20104 1221 20146
rect 1255 20104 1297 20146
rect 1177 20074 1297 20104
rect 1177 20036 1221 20074
rect 1255 20036 1297 20074
rect 1177 20002 1297 20036
rect 1177 19968 1221 20002
rect 1255 19968 1297 20002
rect 1177 19934 1297 19968
rect 1177 19896 1221 19934
rect 1255 19896 1297 19934
rect 1177 19866 1297 19896
rect 1177 19824 1221 19866
rect 1255 19824 1297 19866
rect 1177 19798 1297 19824
rect 1177 19752 1221 19798
rect 1255 19752 1297 19798
rect 1177 19730 1297 19752
rect 1177 19680 1221 19730
rect 1255 19680 1297 19730
rect 1177 19662 1297 19680
rect 1177 19608 1221 19662
rect 1255 19608 1297 19662
rect 1177 19594 1297 19608
rect 1177 19536 1221 19594
rect 1255 19536 1297 19594
rect 1177 19526 1297 19536
rect 1177 19464 1221 19526
rect 1255 19464 1297 19526
rect 1177 19458 1297 19464
rect 1177 19392 1221 19458
rect 1255 19392 1297 19458
rect 1177 19390 1297 19392
rect 1177 19356 1221 19390
rect 1255 19356 1297 19390
rect 1177 19354 1297 19356
rect 1177 19288 1221 19354
rect 1255 19288 1297 19354
rect 1177 19282 1297 19288
rect 1177 19220 1221 19282
rect 1255 19220 1297 19282
rect 1177 19210 1297 19220
rect 1177 19152 1221 19210
rect 1255 19152 1297 19210
rect 1177 19138 1297 19152
rect 1177 19084 1221 19138
rect 1255 19084 1297 19138
rect 1177 19066 1297 19084
rect 1177 19016 1221 19066
rect 1255 19016 1297 19066
rect 1177 18994 1297 19016
rect 1177 18948 1221 18994
rect 1255 18948 1297 18994
rect 1177 18922 1297 18948
rect 1177 18880 1221 18922
rect 1255 18880 1297 18922
rect 1177 18850 1297 18880
rect 1177 18812 1221 18850
rect 1255 18812 1297 18850
rect 1177 18778 1297 18812
rect 1177 18744 1221 18778
rect 1255 18744 1297 18778
rect 1177 18710 1297 18744
rect 1177 18672 1221 18710
rect 1255 18672 1297 18710
rect 1177 18642 1297 18672
rect 1177 18600 1221 18642
rect 1255 18600 1297 18642
rect 1177 18574 1297 18600
rect 1177 18528 1221 18574
rect 1255 18528 1297 18574
rect 1177 18506 1297 18528
rect 1177 18456 1221 18506
rect 1255 18456 1297 18506
rect 1177 18438 1297 18456
rect 1177 18384 1221 18438
rect 1255 18384 1297 18438
rect 1177 18370 1297 18384
rect 1177 18312 1221 18370
rect 1255 18312 1297 18370
rect 1177 18302 1297 18312
rect 1177 18240 1221 18302
rect 1255 18240 1297 18302
rect 1177 18234 1297 18240
rect 1177 18168 1221 18234
rect 1255 18168 1297 18234
rect 1177 18166 1297 18168
rect 1177 18132 1221 18166
rect 1255 18132 1297 18166
rect 1177 18130 1297 18132
rect 1177 18064 1221 18130
rect 1255 18064 1297 18130
rect 1177 18058 1297 18064
rect 1177 17996 1221 18058
rect 1255 17996 1297 18058
rect 1177 17986 1297 17996
rect 1177 17928 1221 17986
rect 1255 17928 1297 17986
rect 1177 17914 1297 17928
rect 1177 17860 1221 17914
rect 1255 17860 1297 17914
rect 1177 17842 1297 17860
rect 1177 17792 1221 17842
rect 1255 17792 1297 17842
rect 1177 17770 1297 17792
rect 1177 17724 1221 17770
rect 1255 17724 1297 17770
rect 1177 17698 1297 17724
rect 1177 17656 1221 17698
rect 1255 17656 1297 17698
rect 1177 17626 1297 17656
rect 1177 17588 1221 17626
rect 1255 17588 1297 17626
rect 1177 17554 1297 17588
rect 1177 17520 1221 17554
rect 1255 17520 1297 17554
rect 1177 17486 1297 17520
rect 1177 17448 1221 17486
rect 1255 17448 1297 17486
rect 1177 17418 1297 17448
rect 1177 17376 1221 17418
rect 1255 17376 1297 17418
rect 1177 17350 1297 17376
rect 1177 17304 1221 17350
rect 1255 17304 1297 17350
rect 1177 17282 1297 17304
rect 1177 17232 1221 17282
rect 1255 17232 1297 17282
rect 1177 17214 1297 17232
rect 1177 17160 1221 17214
rect 1255 17160 1297 17214
rect 1177 17146 1297 17160
rect 1177 17088 1221 17146
rect 1255 17088 1297 17146
rect 1177 17078 1297 17088
rect 1177 17016 1221 17078
rect 1255 17016 1297 17078
rect 1177 17010 1297 17016
rect 1177 16944 1221 17010
rect 1255 16944 1297 17010
rect 1177 16942 1297 16944
rect 1177 16908 1221 16942
rect 1255 16908 1297 16942
rect 1177 16906 1297 16908
rect 1177 16840 1221 16906
rect 1255 16840 1297 16906
rect 1177 16834 1297 16840
rect 1177 16772 1221 16834
rect 1255 16772 1297 16834
rect 1177 16762 1297 16772
rect 1177 16704 1221 16762
rect 1255 16704 1297 16762
rect 1177 16690 1297 16704
rect 1177 16636 1221 16690
rect 1255 16636 1297 16690
rect 1177 16618 1297 16636
rect 1177 16568 1221 16618
rect 1255 16568 1297 16618
rect 1177 16546 1297 16568
rect 1177 16500 1221 16546
rect 1255 16500 1297 16546
rect 1177 16474 1297 16500
rect 1177 16432 1221 16474
rect 1255 16432 1297 16474
rect 1177 16402 1297 16432
rect 1177 16364 1221 16402
rect 1255 16364 1297 16402
rect 1177 16330 1297 16364
rect 1177 16296 1221 16330
rect 1255 16296 1297 16330
rect 1177 16262 1297 16296
rect 1177 16224 1221 16262
rect 1255 16224 1297 16262
rect 1177 16194 1297 16224
rect 1177 16152 1221 16194
rect 1255 16152 1297 16194
rect 1177 16126 1297 16152
rect 1177 16080 1221 16126
rect 1255 16080 1297 16126
rect 1177 16058 1297 16080
rect 1177 16008 1221 16058
rect 1255 16008 1297 16058
rect 1177 15990 1297 16008
rect 1177 15936 1221 15990
rect 1255 15936 1297 15990
rect 1177 15922 1297 15936
rect 1177 15864 1221 15922
rect 1255 15864 1297 15922
rect 1177 15854 1297 15864
rect 1177 15792 1221 15854
rect 1255 15792 1297 15854
rect 1177 15786 1297 15792
rect 1177 15720 1221 15786
rect 1255 15720 1297 15786
rect 1177 15718 1297 15720
rect 1177 15684 1221 15718
rect 1255 15684 1297 15718
rect 1177 15682 1297 15684
rect 1177 15616 1221 15682
rect 1255 15616 1297 15682
rect 1177 15610 1297 15616
rect 1177 15548 1221 15610
rect 1255 15548 1297 15610
rect 1177 15538 1297 15548
rect 1177 15480 1221 15538
rect 1255 15480 1297 15538
rect 1177 15466 1297 15480
rect 1177 15412 1221 15466
rect 1255 15412 1297 15466
rect 1177 15394 1297 15412
rect 1177 15344 1221 15394
rect 1255 15344 1297 15394
rect 1177 15322 1297 15344
rect 1177 15276 1221 15322
rect 1255 15276 1297 15322
rect 1177 15250 1297 15276
rect 1177 15208 1221 15250
rect 1255 15208 1297 15250
rect 1177 15178 1297 15208
rect 1177 15140 1221 15178
rect 1255 15140 1297 15178
rect 1177 15106 1297 15140
rect 1177 15072 1221 15106
rect 1255 15072 1297 15106
rect 1177 15038 1297 15072
rect 1177 15000 1221 15038
rect 1255 15000 1297 15038
rect 1177 14970 1297 15000
rect 1177 14928 1221 14970
rect 1255 14928 1297 14970
rect 1177 14902 1297 14928
rect 1177 14856 1221 14902
rect 1255 14856 1297 14902
rect 1177 14834 1297 14856
rect 1177 14784 1221 14834
rect 1255 14784 1297 14834
rect 1177 14766 1297 14784
rect 1177 14712 1221 14766
rect 1255 14712 1297 14766
rect 1177 14698 1297 14712
rect 1177 14640 1221 14698
rect 1255 14640 1297 14698
rect 1177 14630 1297 14640
rect 1177 14568 1221 14630
rect 1255 14568 1297 14630
rect 1177 14562 1297 14568
rect 1177 14496 1221 14562
rect 1255 14496 1297 14562
rect 1177 14494 1297 14496
rect 1177 14460 1221 14494
rect 1255 14460 1297 14494
rect 1177 14458 1297 14460
rect 1177 14392 1221 14458
rect 1255 14392 1297 14458
rect 1177 14386 1297 14392
rect 1177 14324 1221 14386
rect 1255 14324 1297 14386
rect 1177 14314 1297 14324
rect 1177 14256 1221 14314
rect 1255 14256 1297 14314
rect 1177 14242 1297 14256
rect 1177 14188 1221 14242
rect 1255 14188 1297 14242
rect 1177 14170 1297 14188
rect 1177 14120 1221 14170
rect 1255 14120 1297 14170
rect 1177 14098 1297 14120
rect 1177 14052 1221 14098
rect 1255 14052 1297 14098
rect 1177 14026 1297 14052
rect 1177 13984 1221 14026
rect 1255 13984 1297 14026
rect 1177 13954 1297 13984
rect 1177 13916 1221 13954
rect 1255 13916 1297 13954
rect 1177 13882 1297 13916
rect 1177 13848 1221 13882
rect 1255 13848 1297 13882
rect 1177 13814 1297 13848
rect 1177 13776 1221 13814
rect 1255 13776 1297 13814
rect 1177 13746 1297 13776
rect 1177 13704 1221 13746
rect 1255 13704 1297 13746
rect 1177 13678 1297 13704
rect 1177 13632 1221 13678
rect 1255 13632 1297 13678
rect 1177 13610 1297 13632
rect 1177 13560 1221 13610
rect 1255 13560 1297 13610
rect 1177 13542 1297 13560
rect 1177 13488 1221 13542
rect 1255 13488 1297 13542
rect 1177 13474 1297 13488
rect 1177 13416 1221 13474
rect 1255 13416 1297 13474
rect 1177 13406 1297 13416
rect 1177 13344 1221 13406
rect 1255 13344 1297 13406
rect 1177 13338 1297 13344
rect 1177 13272 1221 13338
rect 1255 13272 1297 13338
rect 1177 13270 1297 13272
rect 1177 13236 1221 13270
rect 1255 13236 1297 13270
rect 1177 13234 1297 13236
rect 1177 13168 1221 13234
rect 1255 13168 1297 13234
rect 1177 13162 1297 13168
rect 1177 13100 1221 13162
rect 1255 13100 1297 13162
rect 1177 13090 1297 13100
rect 1177 13032 1221 13090
rect 1255 13032 1297 13090
rect 1177 13018 1297 13032
rect 1177 12964 1221 13018
rect 1255 12964 1297 13018
rect 1177 12946 1297 12964
rect 1177 12896 1221 12946
rect 1255 12896 1297 12946
rect 1177 12874 1297 12896
rect 1177 12828 1221 12874
rect 1255 12828 1297 12874
rect 1177 12802 1297 12828
rect 1177 12760 1221 12802
rect 1255 12760 1297 12802
rect 1177 12730 1297 12760
rect 1177 12692 1221 12730
rect 1255 12692 1297 12730
rect 1177 12658 1297 12692
rect 1177 12624 1221 12658
rect 1255 12624 1297 12658
rect 1177 12590 1297 12624
rect 1177 12552 1221 12590
rect 1255 12552 1297 12590
rect 1177 12522 1297 12552
rect 1177 12480 1221 12522
rect 1255 12480 1297 12522
rect 1177 12454 1297 12480
rect 1177 12408 1221 12454
rect 1255 12408 1297 12454
rect 1177 12386 1297 12408
rect 1177 12336 1221 12386
rect 1255 12336 1297 12386
rect 1177 12318 1297 12336
rect 1177 12264 1221 12318
rect 1255 12264 1297 12318
rect 1177 12250 1297 12264
rect 1177 12192 1221 12250
rect 1255 12192 1297 12250
rect 1177 12182 1297 12192
rect 1177 12120 1221 12182
rect 1255 12120 1297 12182
rect 1177 12114 1297 12120
rect 1177 12048 1221 12114
rect 1255 12048 1297 12114
rect 1177 12046 1297 12048
rect 1177 12012 1221 12046
rect 1255 12012 1297 12046
rect 1177 12010 1297 12012
rect 1177 11944 1221 12010
rect 1255 11944 1297 12010
rect 1177 11938 1297 11944
rect 1177 11876 1221 11938
rect 1255 11876 1297 11938
rect 1177 11866 1297 11876
rect 1177 11808 1221 11866
rect 1255 11808 1297 11866
rect 1177 11794 1297 11808
rect 1177 11740 1221 11794
rect 1255 11740 1297 11794
rect 1177 11722 1297 11740
rect 1177 11672 1221 11722
rect 1255 11672 1297 11722
rect 1177 11650 1297 11672
rect 1177 11604 1221 11650
rect 1255 11604 1297 11650
rect 1177 11578 1297 11604
rect 1177 11536 1221 11578
rect 1255 11536 1297 11578
rect 1177 11506 1297 11536
rect 1177 11468 1221 11506
rect 1255 11468 1297 11506
rect 1177 11434 1297 11468
rect 1177 11400 1221 11434
rect 1255 11400 1297 11434
rect 1177 11366 1297 11400
rect 1177 11328 1221 11366
rect 1255 11328 1297 11366
rect 1177 11298 1297 11328
rect 1177 11256 1221 11298
rect 1255 11256 1297 11298
rect 1177 11230 1297 11256
rect 1177 11184 1221 11230
rect 1255 11184 1297 11230
rect 1177 11162 1297 11184
rect 1177 11112 1221 11162
rect 1255 11112 1297 11162
rect 1177 11094 1297 11112
rect 1177 11040 1221 11094
rect 1255 11040 1297 11094
rect 1177 11026 1297 11040
rect 1177 10968 1221 11026
rect 1255 10968 1297 11026
rect 1177 10958 1297 10968
rect 1177 10896 1221 10958
rect 1255 10896 1297 10958
rect 1177 10890 1297 10896
rect 1177 10824 1221 10890
rect 1255 10824 1297 10890
rect 1177 10822 1297 10824
rect 1177 10788 1221 10822
rect 1255 10788 1297 10822
rect 1177 10786 1297 10788
rect 1177 10720 1221 10786
rect 1255 10720 1297 10786
rect 1177 10714 1297 10720
rect 1177 10652 1221 10714
rect 1255 10652 1297 10714
rect 1177 10642 1297 10652
rect 1177 10584 1221 10642
rect 1255 10584 1297 10642
rect 1177 10570 1297 10584
rect 1177 10516 1221 10570
rect 1255 10516 1297 10570
rect 1177 10498 1297 10516
rect 1177 10448 1221 10498
rect 1255 10448 1297 10498
rect 1177 10426 1297 10448
rect 1177 10380 1221 10426
rect 1255 10380 1297 10426
rect 1177 10334 1297 10380
rect 13697 34490 13817 34564
rect 13697 34444 13739 34490
rect 13773 34444 13817 34490
rect 13697 34422 13817 34444
rect 13697 34372 13739 34422
rect 13773 34372 13817 34422
rect 13697 34354 13817 34372
rect 13697 34300 13739 34354
rect 13773 34300 13817 34354
rect 13697 34286 13817 34300
rect 13697 34228 13739 34286
rect 13773 34228 13817 34286
rect 13697 34218 13817 34228
rect 13697 34156 13739 34218
rect 13773 34156 13817 34218
rect 13697 34150 13817 34156
rect 13697 34084 13739 34150
rect 13773 34084 13817 34150
rect 13697 34082 13817 34084
rect 13697 34048 13739 34082
rect 13773 34048 13817 34082
rect 13697 34046 13817 34048
rect 13697 33980 13739 34046
rect 13773 33980 13817 34046
rect 13697 33974 13817 33980
rect 13697 33912 13739 33974
rect 13773 33912 13817 33974
rect 13697 33902 13817 33912
rect 13697 33844 13739 33902
rect 13773 33844 13817 33902
rect 13697 33830 13817 33844
rect 13697 33776 13739 33830
rect 13773 33776 13817 33830
rect 13697 33758 13817 33776
rect 13697 33708 13739 33758
rect 13773 33708 13817 33758
rect 13697 33686 13817 33708
rect 13697 33640 13739 33686
rect 13773 33640 13817 33686
rect 13697 33614 13817 33640
rect 13697 33572 13739 33614
rect 13773 33572 13817 33614
rect 13697 33542 13817 33572
rect 13697 33504 13739 33542
rect 13773 33504 13817 33542
rect 13697 33470 13817 33504
rect 13697 33436 13739 33470
rect 13773 33436 13817 33470
rect 13697 33402 13817 33436
rect 13697 33364 13739 33402
rect 13773 33364 13817 33402
rect 13697 33334 13817 33364
rect 13697 33292 13739 33334
rect 13773 33292 13817 33334
rect 13697 33266 13817 33292
rect 13697 33220 13739 33266
rect 13773 33220 13817 33266
rect 13697 33198 13817 33220
rect 13697 33148 13739 33198
rect 13773 33148 13817 33198
rect 13697 33130 13817 33148
rect 13697 33076 13739 33130
rect 13773 33076 13817 33130
rect 13697 33062 13817 33076
rect 13697 33004 13739 33062
rect 13773 33004 13817 33062
rect 13697 32994 13817 33004
rect 13697 32932 13739 32994
rect 13773 32932 13817 32994
rect 13697 32926 13817 32932
rect 13697 32860 13739 32926
rect 13773 32860 13817 32926
rect 13697 32858 13817 32860
rect 13697 32824 13739 32858
rect 13773 32824 13817 32858
rect 13697 32822 13817 32824
rect 13697 32756 13739 32822
rect 13773 32756 13817 32822
rect 13697 32750 13817 32756
rect 13697 32688 13739 32750
rect 13773 32688 13817 32750
rect 13697 32678 13817 32688
rect 13697 32620 13739 32678
rect 13773 32620 13817 32678
rect 13697 32606 13817 32620
rect 13697 32552 13739 32606
rect 13773 32552 13817 32606
rect 13697 32534 13817 32552
rect 13697 32484 13739 32534
rect 13773 32484 13817 32534
rect 13697 32462 13817 32484
rect 13697 32416 13739 32462
rect 13773 32416 13817 32462
rect 13697 32390 13817 32416
rect 13697 32348 13739 32390
rect 13773 32348 13817 32390
rect 13697 32318 13817 32348
rect 13697 32280 13739 32318
rect 13773 32280 13817 32318
rect 13697 32246 13817 32280
rect 13697 32212 13739 32246
rect 13773 32212 13817 32246
rect 13697 32178 13817 32212
rect 13697 32140 13739 32178
rect 13773 32140 13817 32178
rect 13697 32110 13817 32140
rect 13697 32068 13739 32110
rect 13773 32068 13817 32110
rect 13697 32042 13817 32068
rect 13697 31996 13739 32042
rect 13773 31996 13817 32042
rect 13697 31974 13817 31996
rect 13697 31924 13739 31974
rect 13773 31924 13817 31974
rect 13697 31906 13817 31924
rect 13697 31852 13739 31906
rect 13773 31852 13817 31906
rect 13697 31838 13817 31852
rect 13697 31780 13739 31838
rect 13773 31780 13817 31838
rect 13697 31770 13817 31780
rect 13697 31708 13739 31770
rect 13773 31708 13817 31770
rect 13697 31702 13817 31708
rect 13697 31636 13739 31702
rect 13773 31636 13817 31702
rect 13697 31634 13817 31636
rect 13697 31600 13739 31634
rect 13773 31600 13817 31634
rect 13697 31598 13817 31600
rect 13697 31532 13739 31598
rect 13773 31532 13817 31598
rect 13697 31526 13817 31532
rect 13697 31464 13739 31526
rect 13773 31464 13817 31526
rect 13697 31454 13817 31464
rect 13697 31396 13739 31454
rect 13773 31396 13817 31454
rect 13697 31382 13817 31396
rect 13697 31328 13739 31382
rect 13773 31328 13817 31382
rect 13697 31310 13817 31328
rect 13697 31260 13739 31310
rect 13773 31260 13817 31310
rect 13697 31238 13817 31260
rect 13697 31192 13739 31238
rect 13773 31192 13817 31238
rect 13697 31166 13817 31192
rect 13697 31124 13739 31166
rect 13773 31124 13817 31166
rect 13697 31094 13817 31124
rect 13697 31056 13739 31094
rect 13773 31056 13817 31094
rect 13697 31022 13817 31056
rect 13697 30988 13739 31022
rect 13773 30988 13817 31022
rect 13697 30954 13817 30988
rect 13697 30916 13739 30954
rect 13773 30916 13817 30954
rect 13697 30886 13817 30916
rect 13697 30844 13739 30886
rect 13773 30844 13817 30886
rect 13697 30818 13817 30844
rect 13697 30772 13739 30818
rect 13773 30772 13817 30818
rect 13697 30750 13817 30772
rect 13697 30700 13739 30750
rect 13773 30700 13817 30750
rect 13697 30682 13817 30700
rect 13697 30628 13739 30682
rect 13773 30628 13817 30682
rect 13697 30614 13817 30628
rect 13697 30556 13739 30614
rect 13773 30556 13817 30614
rect 13697 30546 13817 30556
rect 13697 30484 13739 30546
rect 13773 30484 13817 30546
rect 13697 30478 13817 30484
rect 13697 30412 13739 30478
rect 13773 30412 13817 30478
rect 13697 30410 13817 30412
rect 13697 30376 13739 30410
rect 13773 30376 13817 30410
rect 13697 30374 13817 30376
rect 13697 30308 13739 30374
rect 13773 30308 13817 30374
rect 13697 30302 13817 30308
rect 13697 30240 13739 30302
rect 13773 30240 13817 30302
rect 13697 30230 13817 30240
rect 13697 30172 13739 30230
rect 13773 30172 13817 30230
rect 13697 30158 13817 30172
rect 13697 30104 13739 30158
rect 13773 30104 13817 30158
rect 13697 30086 13817 30104
rect 13697 30036 13739 30086
rect 13773 30036 13817 30086
rect 13697 30014 13817 30036
rect 13697 29968 13739 30014
rect 13773 29968 13817 30014
rect 13697 29942 13817 29968
rect 13697 29900 13739 29942
rect 13773 29900 13817 29942
rect 13697 29870 13817 29900
rect 13697 29832 13739 29870
rect 13773 29832 13817 29870
rect 13697 29798 13817 29832
rect 13697 29764 13739 29798
rect 13773 29764 13817 29798
rect 13697 29730 13817 29764
rect 13697 29692 13739 29730
rect 13773 29692 13817 29730
rect 13697 29662 13817 29692
rect 13697 29620 13739 29662
rect 13773 29620 13817 29662
rect 13697 29594 13817 29620
rect 13697 29548 13739 29594
rect 13773 29548 13817 29594
rect 13697 29526 13817 29548
rect 13697 29476 13739 29526
rect 13773 29476 13817 29526
rect 13697 29458 13817 29476
rect 13697 29404 13739 29458
rect 13773 29404 13817 29458
rect 13697 29390 13817 29404
rect 13697 29332 13739 29390
rect 13773 29332 13817 29390
rect 13697 29322 13817 29332
rect 13697 29260 13739 29322
rect 13773 29260 13817 29322
rect 13697 29254 13817 29260
rect 13697 29188 13739 29254
rect 13773 29188 13817 29254
rect 13697 29186 13817 29188
rect 13697 29152 13739 29186
rect 13773 29152 13817 29186
rect 13697 29150 13817 29152
rect 13697 29084 13739 29150
rect 13773 29084 13817 29150
rect 13697 29078 13817 29084
rect 13697 29016 13739 29078
rect 13773 29016 13817 29078
rect 13697 29006 13817 29016
rect 13697 28948 13739 29006
rect 13773 28948 13817 29006
rect 13697 28934 13817 28948
rect 13697 28880 13739 28934
rect 13773 28880 13817 28934
rect 13697 28862 13817 28880
rect 13697 28812 13739 28862
rect 13773 28812 13817 28862
rect 13697 28790 13817 28812
rect 13697 28744 13739 28790
rect 13773 28744 13817 28790
rect 13697 28718 13817 28744
rect 13697 28676 13739 28718
rect 13773 28676 13817 28718
rect 13697 28646 13817 28676
rect 13697 28608 13739 28646
rect 13773 28608 13817 28646
rect 13697 28574 13817 28608
rect 13697 28540 13739 28574
rect 13773 28540 13817 28574
rect 13697 28506 13817 28540
rect 13697 28468 13739 28506
rect 13773 28468 13817 28506
rect 13697 28438 13817 28468
rect 13697 28396 13739 28438
rect 13773 28396 13817 28438
rect 13697 28370 13817 28396
rect 13697 28324 13739 28370
rect 13773 28324 13817 28370
rect 13697 28302 13817 28324
rect 13697 28252 13739 28302
rect 13773 28252 13817 28302
rect 13697 28234 13817 28252
rect 13697 28180 13739 28234
rect 13773 28180 13817 28234
rect 13697 28166 13817 28180
rect 13697 28108 13739 28166
rect 13773 28108 13817 28166
rect 13697 28098 13817 28108
rect 13697 28036 13739 28098
rect 13773 28036 13817 28098
rect 13697 28030 13817 28036
rect 13697 27964 13739 28030
rect 13773 27964 13817 28030
rect 13697 27962 13817 27964
rect 13697 27928 13739 27962
rect 13773 27928 13817 27962
rect 13697 27926 13817 27928
rect 13697 27860 13739 27926
rect 13773 27860 13817 27926
rect 13697 27854 13817 27860
rect 13697 27792 13739 27854
rect 13773 27792 13817 27854
rect 13697 27782 13817 27792
rect 13697 27724 13739 27782
rect 13773 27724 13817 27782
rect 13697 27710 13817 27724
rect 13697 27656 13739 27710
rect 13773 27656 13817 27710
rect 13697 27638 13817 27656
rect 13697 27588 13739 27638
rect 13773 27588 13817 27638
rect 13697 27566 13817 27588
rect 13697 27520 13739 27566
rect 13773 27520 13817 27566
rect 13697 27494 13817 27520
rect 13697 27452 13739 27494
rect 13773 27452 13817 27494
rect 13697 27422 13817 27452
rect 13697 27384 13739 27422
rect 13773 27384 13817 27422
rect 13697 27350 13817 27384
rect 13697 27316 13739 27350
rect 13773 27316 13817 27350
rect 13697 27282 13817 27316
rect 13697 27244 13739 27282
rect 13773 27244 13817 27282
rect 13697 27214 13817 27244
rect 13697 27172 13739 27214
rect 13773 27172 13817 27214
rect 13697 27146 13817 27172
rect 13697 27100 13739 27146
rect 13773 27100 13817 27146
rect 13697 27078 13817 27100
rect 13697 27028 13739 27078
rect 13773 27028 13817 27078
rect 13697 27010 13817 27028
rect 13697 26956 13739 27010
rect 13773 26956 13817 27010
rect 13697 26942 13817 26956
rect 13697 26884 13739 26942
rect 13773 26884 13817 26942
rect 13697 26874 13817 26884
rect 13697 26812 13739 26874
rect 13773 26812 13817 26874
rect 13697 26806 13817 26812
rect 13697 26740 13739 26806
rect 13773 26740 13817 26806
rect 13697 26738 13817 26740
rect 13697 26704 13739 26738
rect 13773 26704 13817 26738
rect 13697 26702 13817 26704
rect 13697 26636 13739 26702
rect 13773 26636 13817 26702
rect 13697 26630 13817 26636
rect 13697 26568 13739 26630
rect 13773 26568 13817 26630
rect 13697 26558 13817 26568
rect 13697 26500 13739 26558
rect 13773 26500 13817 26558
rect 13697 26486 13817 26500
rect 13697 26432 13739 26486
rect 13773 26432 13817 26486
rect 13697 26414 13817 26432
rect 13697 26364 13739 26414
rect 13773 26364 13817 26414
rect 13697 26342 13817 26364
rect 13697 26296 13739 26342
rect 13773 26296 13817 26342
rect 13697 26270 13817 26296
rect 13697 26228 13739 26270
rect 13773 26228 13817 26270
rect 13697 26198 13817 26228
rect 13697 26160 13739 26198
rect 13773 26160 13817 26198
rect 13697 26126 13817 26160
rect 13697 26092 13739 26126
rect 13773 26092 13817 26126
rect 13697 26058 13817 26092
rect 13697 26020 13739 26058
rect 13773 26020 13817 26058
rect 13697 25990 13817 26020
rect 13697 25948 13739 25990
rect 13773 25948 13817 25990
rect 13697 25922 13817 25948
rect 13697 25876 13739 25922
rect 13773 25876 13817 25922
rect 13697 25854 13817 25876
rect 13697 25804 13739 25854
rect 13773 25804 13817 25854
rect 13697 25786 13817 25804
rect 13697 25732 13739 25786
rect 13773 25732 13817 25786
rect 13697 25718 13817 25732
rect 13697 25660 13739 25718
rect 13773 25660 13817 25718
rect 13697 25650 13817 25660
rect 13697 25588 13739 25650
rect 13773 25588 13817 25650
rect 13697 25582 13817 25588
rect 13697 25516 13739 25582
rect 13773 25516 13817 25582
rect 13697 25514 13817 25516
rect 13697 25480 13739 25514
rect 13773 25480 13817 25514
rect 13697 25478 13817 25480
rect 13697 25412 13739 25478
rect 13773 25412 13817 25478
rect 13697 25406 13817 25412
rect 13697 25344 13739 25406
rect 13773 25344 13817 25406
rect 13697 25334 13817 25344
rect 13697 25276 13739 25334
rect 13773 25276 13817 25334
rect 13697 25262 13817 25276
rect 13697 25208 13739 25262
rect 13773 25208 13817 25262
rect 13697 25190 13817 25208
rect 13697 25140 13739 25190
rect 13773 25140 13817 25190
rect 13697 25118 13817 25140
rect 13697 25072 13739 25118
rect 13773 25072 13817 25118
rect 13697 25046 13817 25072
rect 13697 25004 13739 25046
rect 13773 25004 13817 25046
rect 13697 24974 13817 25004
rect 13697 24936 13739 24974
rect 13773 24936 13817 24974
rect 13697 24902 13817 24936
rect 13697 24868 13739 24902
rect 13773 24868 13817 24902
rect 13697 24834 13817 24868
rect 13697 24796 13739 24834
rect 13773 24796 13817 24834
rect 13697 24766 13817 24796
rect 13697 24724 13739 24766
rect 13773 24724 13817 24766
rect 13697 24698 13817 24724
rect 13697 24652 13739 24698
rect 13773 24652 13817 24698
rect 13697 24630 13817 24652
rect 13697 24580 13739 24630
rect 13773 24580 13817 24630
rect 13697 24562 13817 24580
rect 13697 24508 13739 24562
rect 13773 24508 13817 24562
rect 13697 24494 13817 24508
rect 13697 24436 13739 24494
rect 13773 24436 13817 24494
rect 13697 24426 13817 24436
rect 13697 24364 13739 24426
rect 13773 24364 13817 24426
rect 13697 24358 13817 24364
rect 13697 24292 13739 24358
rect 13773 24292 13817 24358
rect 13697 24290 13817 24292
rect 13697 24256 13739 24290
rect 13773 24256 13817 24290
rect 13697 24254 13817 24256
rect 13697 24188 13739 24254
rect 13773 24188 13817 24254
rect 13697 24182 13817 24188
rect 13697 24120 13739 24182
rect 13773 24120 13817 24182
rect 13697 24110 13817 24120
rect 13697 24052 13739 24110
rect 13773 24052 13817 24110
rect 13697 24038 13817 24052
rect 13697 23984 13739 24038
rect 13773 23984 13817 24038
rect 13697 23966 13817 23984
rect 13697 23916 13739 23966
rect 13773 23916 13817 23966
rect 13697 23894 13817 23916
rect 13697 23848 13739 23894
rect 13773 23848 13817 23894
rect 13697 23822 13817 23848
rect 13697 23780 13739 23822
rect 13773 23780 13817 23822
rect 13697 23750 13817 23780
rect 13697 23712 13739 23750
rect 13773 23712 13817 23750
rect 13697 23678 13817 23712
rect 13697 23644 13739 23678
rect 13773 23644 13817 23678
rect 13697 23610 13817 23644
rect 13697 23572 13739 23610
rect 13773 23572 13817 23610
rect 13697 23542 13817 23572
rect 13697 23500 13739 23542
rect 13773 23500 13817 23542
rect 13697 23474 13817 23500
rect 13697 23428 13739 23474
rect 13773 23428 13817 23474
rect 13697 23406 13817 23428
rect 13697 23356 13739 23406
rect 13773 23356 13817 23406
rect 13697 23338 13817 23356
rect 13697 23284 13739 23338
rect 13773 23284 13817 23338
rect 13697 23270 13817 23284
rect 13697 23212 13739 23270
rect 13773 23212 13817 23270
rect 13697 23202 13817 23212
rect 13697 23140 13739 23202
rect 13773 23140 13817 23202
rect 13697 23134 13817 23140
rect 13697 23068 13739 23134
rect 13773 23068 13817 23134
rect 13697 23066 13817 23068
rect 13697 23032 13739 23066
rect 13773 23032 13817 23066
rect 13697 23030 13817 23032
rect 13697 22964 13739 23030
rect 13773 22964 13817 23030
rect 13697 22958 13817 22964
rect 13697 22896 13739 22958
rect 13773 22896 13817 22958
rect 13697 22886 13817 22896
rect 13697 22828 13739 22886
rect 13773 22828 13817 22886
rect 13697 22814 13817 22828
rect 13697 22760 13739 22814
rect 13773 22760 13817 22814
rect 13697 22742 13817 22760
rect 13697 22692 13739 22742
rect 13773 22692 13817 22742
rect 13697 22670 13817 22692
rect 13697 22624 13739 22670
rect 13773 22624 13817 22670
rect 13697 22598 13817 22624
rect 13697 22556 13739 22598
rect 13773 22556 13817 22598
rect 13697 22526 13817 22556
rect 13697 22488 13739 22526
rect 13773 22488 13817 22526
rect 13697 22454 13817 22488
rect 13697 22420 13739 22454
rect 13773 22420 13817 22454
rect 13697 22386 13817 22420
rect 13697 22348 13739 22386
rect 13773 22348 13817 22386
rect 13697 22318 13817 22348
rect 13697 22276 13739 22318
rect 13773 22276 13817 22318
rect 13697 22250 13817 22276
rect 13697 22204 13739 22250
rect 13773 22204 13817 22250
rect 13697 22182 13817 22204
rect 13697 22132 13739 22182
rect 13773 22132 13817 22182
rect 13697 22114 13817 22132
rect 13697 22060 13739 22114
rect 13773 22060 13817 22114
rect 13697 22046 13817 22060
rect 13697 21988 13739 22046
rect 13773 21988 13817 22046
rect 13697 21978 13817 21988
rect 13697 21916 13739 21978
rect 13773 21916 13817 21978
rect 13697 21910 13817 21916
rect 13697 21844 13739 21910
rect 13773 21844 13817 21910
rect 13697 21842 13817 21844
rect 13697 21808 13739 21842
rect 13773 21808 13817 21842
rect 13697 21806 13817 21808
rect 13697 21740 13739 21806
rect 13773 21740 13817 21806
rect 13697 21734 13817 21740
rect 13697 21672 13739 21734
rect 13773 21672 13817 21734
rect 13697 21662 13817 21672
rect 13697 21604 13739 21662
rect 13773 21604 13817 21662
rect 13697 21590 13817 21604
rect 13697 21536 13739 21590
rect 13773 21536 13817 21590
rect 13697 21518 13817 21536
rect 13697 21468 13739 21518
rect 13773 21468 13817 21518
rect 13697 21446 13817 21468
rect 13697 21400 13739 21446
rect 13773 21400 13817 21446
rect 13697 21374 13817 21400
rect 13697 21332 13739 21374
rect 13773 21332 13817 21374
rect 13697 21302 13817 21332
rect 13697 21264 13739 21302
rect 13773 21264 13817 21302
rect 13697 21230 13817 21264
rect 13697 21196 13739 21230
rect 13773 21196 13817 21230
rect 13697 21162 13817 21196
rect 13697 21124 13739 21162
rect 13773 21124 13817 21162
rect 13697 21094 13817 21124
rect 13697 21052 13739 21094
rect 13773 21052 13817 21094
rect 13697 21026 13817 21052
rect 13697 20980 13739 21026
rect 13773 20980 13817 21026
rect 13697 20958 13817 20980
rect 13697 20908 13739 20958
rect 13773 20908 13817 20958
rect 13697 20890 13817 20908
rect 13697 20836 13739 20890
rect 13773 20836 13817 20890
rect 13697 20822 13817 20836
rect 13697 20764 13739 20822
rect 13773 20764 13817 20822
rect 13697 20754 13817 20764
rect 13697 20692 13739 20754
rect 13773 20692 13817 20754
rect 13697 20686 13817 20692
rect 13697 20620 13739 20686
rect 13773 20620 13817 20686
rect 13697 20618 13817 20620
rect 13697 20584 13739 20618
rect 13773 20584 13817 20618
rect 13697 20582 13817 20584
rect 13697 20516 13739 20582
rect 13773 20516 13817 20582
rect 13697 20510 13817 20516
rect 13697 20448 13739 20510
rect 13773 20448 13817 20510
rect 13697 20438 13817 20448
rect 13697 20380 13739 20438
rect 13773 20380 13817 20438
rect 13697 20366 13817 20380
rect 13697 20312 13739 20366
rect 13773 20312 13817 20366
rect 13697 20294 13817 20312
rect 13697 20244 13739 20294
rect 13773 20244 13817 20294
rect 13697 20222 13817 20244
rect 13697 20176 13739 20222
rect 13773 20176 13817 20222
rect 13697 20150 13817 20176
rect 13697 20108 13739 20150
rect 13773 20108 13817 20150
rect 13697 20078 13817 20108
rect 13697 20040 13739 20078
rect 13773 20040 13817 20078
rect 13697 20006 13817 20040
rect 13697 19972 13739 20006
rect 13773 19972 13817 20006
rect 13697 19938 13817 19972
rect 13697 19900 13739 19938
rect 13773 19900 13817 19938
rect 13697 19870 13817 19900
rect 13697 19828 13739 19870
rect 13773 19828 13817 19870
rect 13697 19802 13817 19828
rect 13697 19756 13739 19802
rect 13773 19756 13817 19802
rect 13697 19734 13817 19756
rect 13697 19684 13739 19734
rect 13773 19684 13817 19734
rect 13697 19666 13817 19684
rect 13697 19612 13739 19666
rect 13773 19612 13817 19666
rect 13697 19598 13817 19612
rect 13697 19540 13739 19598
rect 13773 19540 13817 19598
rect 13697 19530 13817 19540
rect 13697 19468 13739 19530
rect 13773 19468 13817 19530
rect 13697 19462 13817 19468
rect 13697 19396 13739 19462
rect 13773 19396 13817 19462
rect 13697 19394 13817 19396
rect 13697 19360 13739 19394
rect 13773 19360 13817 19394
rect 13697 19358 13817 19360
rect 13697 19292 13739 19358
rect 13773 19292 13817 19358
rect 13697 19286 13817 19292
rect 13697 19224 13739 19286
rect 13773 19224 13817 19286
rect 13697 19214 13817 19224
rect 13697 19156 13739 19214
rect 13773 19156 13817 19214
rect 13697 19142 13817 19156
rect 13697 19088 13739 19142
rect 13773 19088 13817 19142
rect 13697 19070 13817 19088
rect 13697 19020 13739 19070
rect 13773 19020 13817 19070
rect 13697 18998 13817 19020
rect 13697 18952 13739 18998
rect 13773 18952 13817 18998
rect 13697 18926 13817 18952
rect 13697 18884 13739 18926
rect 13773 18884 13817 18926
rect 13697 18854 13817 18884
rect 13697 18816 13739 18854
rect 13773 18816 13817 18854
rect 13697 18782 13817 18816
rect 13697 18748 13739 18782
rect 13773 18748 13817 18782
rect 13697 18714 13817 18748
rect 13697 18676 13739 18714
rect 13773 18676 13817 18714
rect 13697 18646 13817 18676
rect 13697 18604 13739 18646
rect 13773 18604 13817 18646
rect 13697 18578 13817 18604
rect 13697 18532 13739 18578
rect 13773 18532 13817 18578
rect 13697 18510 13817 18532
rect 13697 18460 13739 18510
rect 13773 18460 13817 18510
rect 13697 18442 13817 18460
rect 13697 18388 13739 18442
rect 13773 18388 13817 18442
rect 13697 18374 13817 18388
rect 13697 18316 13739 18374
rect 13773 18316 13817 18374
rect 13697 18306 13817 18316
rect 13697 18244 13739 18306
rect 13773 18244 13817 18306
rect 13697 18238 13817 18244
rect 13697 18172 13739 18238
rect 13773 18172 13817 18238
rect 13697 18170 13817 18172
rect 13697 18136 13739 18170
rect 13773 18136 13817 18170
rect 13697 18134 13817 18136
rect 13697 18068 13739 18134
rect 13773 18068 13817 18134
rect 13697 18062 13817 18068
rect 13697 18000 13739 18062
rect 13773 18000 13817 18062
rect 13697 17990 13817 18000
rect 13697 17932 13739 17990
rect 13773 17932 13817 17990
rect 13697 17918 13817 17932
rect 13697 17864 13739 17918
rect 13773 17864 13817 17918
rect 13697 17846 13817 17864
rect 13697 17796 13739 17846
rect 13773 17796 13817 17846
rect 13697 17774 13817 17796
rect 13697 17728 13739 17774
rect 13773 17728 13817 17774
rect 13697 17702 13817 17728
rect 13697 17660 13739 17702
rect 13773 17660 13817 17702
rect 13697 17630 13817 17660
rect 13697 17592 13739 17630
rect 13773 17592 13817 17630
rect 13697 17558 13817 17592
rect 13697 17524 13739 17558
rect 13773 17524 13817 17558
rect 13697 17490 13817 17524
rect 13697 17452 13739 17490
rect 13773 17452 13817 17490
rect 13697 17422 13817 17452
rect 13697 17380 13739 17422
rect 13773 17380 13817 17422
rect 13697 17354 13817 17380
rect 13697 17308 13739 17354
rect 13773 17308 13817 17354
rect 13697 17286 13817 17308
rect 13697 17236 13739 17286
rect 13773 17236 13817 17286
rect 13697 17218 13817 17236
rect 13697 17164 13739 17218
rect 13773 17164 13817 17218
rect 13697 17150 13817 17164
rect 13697 17092 13739 17150
rect 13773 17092 13817 17150
rect 13697 17082 13817 17092
rect 13697 17020 13739 17082
rect 13773 17020 13817 17082
rect 13697 17014 13817 17020
rect 13697 16948 13739 17014
rect 13773 16948 13817 17014
rect 13697 16946 13817 16948
rect 13697 16912 13739 16946
rect 13773 16912 13817 16946
rect 13697 16910 13817 16912
rect 13697 16844 13739 16910
rect 13773 16844 13817 16910
rect 13697 16838 13817 16844
rect 13697 16776 13739 16838
rect 13773 16776 13817 16838
rect 13697 16766 13817 16776
rect 13697 16708 13739 16766
rect 13773 16708 13817 16766
rect 13697 16694 13817 16708
rect 13697 16640 13739 16694
rect 13773 16640 13817 16694
rect 13697 16622 13817 16640
rect 13697 16572 13739 16622
rect 13773 16572 13817 16622
rect 13697 16550 13817 16572
rect 13697 16504 13739 16550
rect 13773 16504 13817 16550
rect 13697 16478 13817 16504
rect 13697 16436 13739 16478
rect 13773 16436 13817 16478
rect 13697 16406 13817 16436
rect 13697 16368 13739 16406
rect 13773 16368 13817 16406
rect 13697 16334 13817 16368
rect 13697 16300 13739 16334
rect 13773 16300 13817 16334
rect 13697 16266 13817 16300
rect 13697 16228 13739 16266
rect 13773 16228 13817 16266
rect 13697 16198 13817 16228
rect 13697 16156 13739 16198
rect 13773 16156 13817 16198
rect 13697 16130 13817 16156
rect 13697 16084 13739 16130
rect 13773 16084 13817 16130
rect 13697 16062 13817 16084
rect 13697 16012 13739 16062
rect 13773 16012 13817 16062
rect 13697 15994 13817 16012
rect 13697 15940 13739 15994
rect 13773 15940 13817 15994
rect 13697 15926 13817 15940
rect 13697 15868 13739 15926
rect 13773 15868 13817 15926
rect 13697 15858 13817 15868
rect 13697 15796 13739 15858
rect 13773 15796 13817 15858
rect 13697 15790 13817 15796
rect 13697 15724 13739 15790
rect 13773 15724 13817 15790
rect 13697 15722 13817 15724
rect 13697 15688 13739 15722
rect 13773 15688 13817 15722
rect 13697 15686 13817 15688
rect 13697 15620 13739 15686
rect 13773 15620 13817 15686
rect 13697 15614 13817 15620
rect 13697 15552 13739 15614
rect 13773 15552 13817 15614
rect 13697 15542 13817 15552
rect 13697 15484 13739 15542
rect 13773 15484 13817 15542
rect 13697 15470 13817 15484
rect 13697 15416 13739 15470
rect 13773 15416 13817 15470
rect 13697 15398 13817 15416
rect 13697 15348 13739 15398
rect 13773 15348 13817 15398
rect 13697 15326 13817 15348
rect 13697 15280 13739 15326
rect 13773 15280 13817 15326
rect 13697 15254 13817 15280
rect 13697 15212 13739 15254
rect 13773 15212 13817 15254
rect 13697 15182 13817 15212
rect 13697 15144 13739 15182
rect 13773 15144 13817 15182
rect 13697 15110 13817 15144
rect 13697 15076 13739 15110
rect 13773 15076 13817 15110
rect 13697 15042 13817 15076
rect 13697 15004 13739 15042
rect 13773 15004 13817 15042
rect 13697 14974 13817 15004
rect 13697 14932 13739 14974
rect 13773 14932 13817 14974
rect 13697 14906 13817 14932
rect 13697 14860 13739 14906
rect 13773 14860 13817 14906
rect 13697 14838 13817 14860
rect 13697 14788 13739 14838
rect 13773 14788 13817 14838
rect 13697 14770 13817 14788
rect 13697 14716 13739 14770
rect 13773 14716 13817 14770
rect 13697 14702 13817 14716
rect 13697 14644 13739 14702
rect 13773 14644 13817 14702
rect 13697 14634 13817 14644
rect 13697 14572 13739 14634
rect 13773 14572 13817 14634
rect 13697 14566 13817 14572
rect 13697 14500 13739 14566
rect 13773 14500 13817 14566
rect 13697 14498 13817 14500
rect 13697 14464 13739 14498
rect 13773 14464 13817 14498
rect 13697 14462 13817 14464
rect 13697 14396 13739 14462
rect 13773 14396 13817 14462
rect 13697 14390 13817 14396
rect 13697 14328 13739 14390
rect 13773 14328 13817 14390
rect 13697 14318 13817 14328
rect 13697 14260 13739 14318
rect 13773 14260 13817 14318
rect 13697 14246 13817 14260
rect 13697 14192 13739 14246
rect 13773 14192 13817 14246
rect 13697 14174 13817 14192
rect 13697 14124 13739 14174
rect 13773 14124 13817 14174
rect 13697 14102 13817 14124
rect 13697 14056 13739 14102
rect 13773 14056 13817 14102
rect 13697 14030 13817 14056
rect 13697 13988 13739 14030
rect 13773 13988 13817 14030
rect 13697 13958 13817 13988
rect 13697 13920 13739 13958
rect 13773 13920 13817 13958
rect 13697 13886 13817 13920
rect 13697 13852 13739 13886
rect 13773 13852 13817 13886
rect 13697 13818 13817 13852
rect 13697 13780 13739 13818
rect 13773 13780 13817 13818
rect 13697 13750 13817 13780
rect 13697 13708 13739 13750
rect 13773 13708 13817 13750
rect 13697 13682 13817 13708
rect 13697 13636 13739 13682
rect 13773 13636 13817 13682
rect 13697 13614 13817 13636
rect 13697 13564 13739 13614
rect 13773 13564 13817 13614
rect 13697 13546 13817 13564
rect 13697 13492 13739 13546
rect 13773 13492 13817 13546
rect 13697 13478 13817 13492
rect 13697 13420 13739 13478
rect 13773 13420 13817 13478
rect 13697 13410 13817 13420
rect 13697 13348 13739 13410
rect 13773 13348 13817 13410
rect 13697 13342 13817 13348
rect 13697 13276 13739 13342
rect 13773 13276 13817 13342
rect 13697 13274 13817 13276
rect 13697 13240 13739 13274
rect 13773 13240 13817 13274
rect 13697 13238 13817 13240
rect 13697 13172 13739 13238
rect 13773 13172 13817 13238
rect 13697 13166 13817 13172
rect 13697 13104 13739 13166
rect 13773 13104 13817 13166
rect 13697 13094 13817 13104
rect 13697 13036 13739 13094
rect 13773 13036 13817 13094
rect 13697 13022 13817 13036
rect 13697 12968 13739 13022
rect 13773 12968 13817 13022
rect 13697 12950 13817 12968
rect 13697 12900 13739 12950
rect 13773 12900 13817 12950
rect 13697 12878 13817 12900
rect 13697 12832 13739 12878
rect 13773 12832 13817 12878
rect 13697 12806 13817 12832
rect 13697 12764 13739 12806
rect 13773 12764 13817 12806
rect 13697 12734 13817 12764
rect 13697 12696 13739 12734
rect 13773 12696 13817 12734
rect 13697 12662 13817 12696
rect 13697 12628 13739 12662
rect 13773 12628 13817 12662
rect 13697 12594 13817 12628
rect 13697 12556 13739 12594
rect 13773 12556 13817 12594
rect 13697 12526 13817 12556
rect 13697 12484 13739 12526
rect 13773 12484 13817 12526
rect 13697 12458 13817 12484
rect 13697 12412 13739 12458
rect 13773 12412 13817 12458
rect 13697 12390 13817 12412
rect 13697 12340 13739 12390
rect 13773 12340 13817 12390
rect 13697 12322 13817 12340
rect 13697 12268 13739 12322
rect 13773 12268 13817 12322
rect 13697 12254 13817 12268
rect 13697 12196 13739 12254
rect 13773 12196 13817 12254
rect 13697 12186 13817 12196
rect 13697 12124 13739 12186
rect 13773 12124 13817 12186
rect 13697 12118 13817 12124
rect 13697 12052 13739 12118
rect 13773 12052 13817 12118
rect 13697 12050 13817 12052
rect 13697 12016 13739 12050
rect 13773 12016 13817 12050
rect 13697 12014 13817 12016
rect 13697 11948 13739 12014
rect 13773 11948 13817 12014
rect 13697 11942 13817 11948
rect 13697 11880 13739 11942
rect 13773 11880 13817 11942
rect 13697 11870 13817 11880
rect 13697 11812 13739 11870
rect 13773 11812 13817 11870
rect 13697 11798 13817 11812
rect 13697 11744 13739 11798
rect 13773 11744 13817 11798
rect 13697 11726 13817 11744
rect 13697 11676 13739 11726
rect 13773 11676 13817 11726
rect 13697 11654 13817 11676
rect 13697 11608 13739 11654
rect 13773 11608 13817 11654
rect 13697 11582 13817 11608
rect 13697 11540 13739 11582
rect 13773 11540 13817 11582
rect 13697 11510 13817 11540
rect 13697 11472 13739 11510
rect 13773 11472 13817 11510
rect 13697 11438 13817 11472
rect 13697 11404 13739 11438
rect 13773 11404 13817 11438
rect 13697 11370 13817 11404
rect 13697 11332 13739 11370
rect 13773 11332 13817 11370
rect 13697 11302 13817 11332
rect 13697 11260 13739 11302
rect 13773 11260 13817 11302
rect 13697 11234 13817 11260
rect 13697 11188 13739 11234
rect 13773 11188 13817 11234
rect 13697 11166 13817 11188
rect 13697 11116 13739 11166
rect 13773 11116 13817 11166
rect 13697 11098 13817 11116
rect 13697 11044 13739 11098
rect 13773 11044 13817 11098
rect 13697 11030 13817 11044
rect 13697 10972 13739 11030
rect 13773 10972 13817 11030
rect 13697 10962 13817 10972
rect 13697 10900 13739 10962
rect 13773 10900 13817 10962
rect 13697 10894 13817 10900
rect 13697 10828 13739 10894
rect 13773 10828 13817 10894
rect 13697 10826 13817 10828
rect 13697 10792 13739 10826
rect 13773 10792 13817 10826
rect 13697 10790 13817 10792
rect 13697 10724 13739 10790
rect 13773 10724 13817 10790
rect 13697 10718 13817 10724
rect 13697 10656 13739 10718
rect 13773 10656 13817 10718
rect 13697 10646 13817 10656
rect 13697 10588 13739 10646
rect 13773 10588 13817 10646
rect 13697 10574 13817 10588
rect 13697 10520 13739 10574
rect 13773 10520 13817 10574
rect 13697 10502 13817 10520
rect 13697 10452 13739 10502
rect 13773 10452 13817 10502
rect 13697 10430 13817 10452
rect 13697 10384 13739 10430
rect 13773 10384 13817 10430
rect 13697 10334 13817 10384
rect 1177 10290 13817 10334
rect 1177 10256 1355 10290
rect 1389 10256 1423 10290
rect 1461 10256 1491 10290
rect 1533 10256 1559 10290
rect 1605 10256 1627 10290
rect 1677 10256 1695 10290
rect 1749 10256 1763 10290
rect 1821 10256 1831 10290
rect 1893 10256 1899 10290
rect 1965 10256 1967 10290
rect 2001 10256 2003 10290
rect 2069 10256 2075 10290
rect 2137 10256 2147 10290
rect 2205 10256 2219 10290
rect 2273 10256 2291 10290
rect 2341 10256 2363 10290
rect 2409 10256 2435 10290
rect 2477 10256 2507 10290
rect 2545 10256 2579 10290
rect 2613 10256 2647 10290
rect 2685 10256 2715 10290
rect 2757 10256 2783 10290
rect 2829 10256 2851 10290
rect 2901 10256 2919 10290
rect 2973 10256 2987 10290
rect 3045 10256 3055 10290
rect 3117 10256 3123 10290
rect 3189 10256 3191 10290
rect 3225 10256 3227 10290
rect 3293 10256 3299 10290
rect 3361 10256 3371 10290
rect 3429 10256 3443 10290
rect 3497 10256 3515 10290
rect 3565 10256 3587 10290
rect 3633 10256 3659 10290
rect 3701 10256 3731 10290
rect 3769 10256 3803 10290
rect 3837 10256 3871 10290
rect 3909 10256 3939 10290
rect 3981 10256 4007 10290
rect 4053 10256 4075 10290
rect 4125 10256 4143 10290
rect 4197 10256 4211 10290
rect 4269 10256 4279 10290
rect 4341 10256 4347 10290
rect 4413 10256 4415 10290
rect 4449 10256 4451 10290
rect 4517 10256 4523 10290
rect 4585 10256 4595 10290
rect 4653 10256 4667 10290
rect 4721 10256 4739 10290
rect 4789 10256 4811 10290
rect 4857 10256 4883 10290
rect 4925 10256 4955 10290
rect 4993 10256 5027 10290
rect 5061 10256 5095 10290
rect 5133 10256 5163 10290
rect 5205 10256 5231 10290
rect 5277 10256 5299 10290
rect 5349 10256 5367 10290
rect 5421 10256 5435 10290
rect 5493 10256 5503 10290
rect 5565 10256 5571 10290
rect 5637 10256 5639 10290
rect 5673 10256 5675 10290
rect 5741 10256 5747 10290
rect 5809 10256 5819 10290
rect 5877 10256 5891 10290
rect 5945 10256 5963 10290
rect 6013 10256 6035 10290
rect 6081 10256 6107 10290
rect 6149 10256 6179 10290
rect 6217 10256 6251 10290
rect 6285 10256 6319 10290
rect 6357 10256 6387 10290
rect 6429 10256 6455 10290
rect 6501 10256 6523 10290
rect 6573 10256 6591 10290
rect 6645 10256 6659 10290
rect 6717 10256 6727 10290
rect 6789 10256 6795 10290
rect 6861 10256 6863 10290
rect 6897 10256 6899 10290
rect 6965 10256 6971 10290
rect 7033 10256 7043 10290
rect 7101 10256 7115 10290
rect 7169 10256 7187 10290
rect 7237 10256 7259 10290
rect 7305 10256 7331 10290
rect 7373 10256 7403 10290
rect 7441 10256 7475 10290
rect 7509 10256 7543 10290
rect 7581 10256 7611 10290
rect 7653 10256 7679 10290
rect 7725 10256 7747 10290
rect 7797 10256 7815 10290
rect 7869 10256 7883 10290
rect 7941 10256 7951 10290
rect 8013 10256 8019 10290
rect 8085 10256 8087 10290
rect 8121 10256 8123 10290
rect 8189 10256 8195 10290
rect 8257 10256 8267 10290
rect 8325 10256 8339 10290
rect 8393 10256 8411 10290
rect 8461 10256 8483 10290
rect 8529 10256 8555 10290
rect 8597 10256 8627 10290
rect 8665 10256 8699 10290
rect 8733 10256 8767 10290
rect 8805 10256 8835 10290
rect 8877 10256 8903 10290
rect 8949 10256 8971 10290
rect 9021 10256 9039 10290
rect 9093 10256 9107 10290
rect 9165 10256 9175 10290
rect 9237 10256 9243 10290
rect 9309 10256 9311 10290
rect 9345 10256 9347 10290
rect 9413 10256 9419 10290
rect 9481 10256 9491 10290
rect 9549 10256 9563 10290
rect 9617 10256 9635 10290
rect 9685 10256 9707 10290
rect 9753 10256 9779 10290
rect 9821 10256 9851 10290
rect 9889 10256 9923 10290
rect 9957 10256 9991 10290
rect 10029 10256 10059 10290
rect 10101 10256 10127 10290
rect 10173 10256 10195 10290
rect 10245 10256 10263 10290
rect 10317 10256 10331 10290
rect 10389 10256 10399 10290
rect 10461 10256 10467 10290
rect 10533 10256 10535 10290
rect 10569 10256 10571 10290
rect 10637 10256 10643 10290
rect 10705 10256 10715 10290
rect 10773 10256 10787 10290
rect 10841 10256 10859 10290
rect 10909 10256 10931 10290
rect 10977 10256 11003 10290
rect 11045 10256 11075 10290
rect 11113 10256 11147 10290
rect 11181 10256 11215 10290
rect 11253 10256 11283 10290
rect 11325 10256 11351 10290
rect 11397 10256 11419 10290
rect 11469 10256 11487 10290
rect 11541 10256 11555 10290
rect 11613 10256 11623 10290
rect 11685 10256 11691 10290
rect 11757 10256 11759 10290
rect 11793 10256 11795 10290
rect 11861 10256 11867 10290
rect 11929 10256 11939 10290
rect 11997 10256 12011 10290
rect 12065 10256 12083 10290
rect 12133 10256 12155 10290
rect 12201 10256 12227 10290
rect 12269 10256 12299 10290
rect 12337 10256 12371 10290
rect 12405 10256 12439 10290
rect 12477 10256 12507 10290
rect 12549 10256 12575 10290
rect 12621 10256 12643 10290
rect 12693 10256 12711 10290
rect 12765 10256 12779 10290
rect 12837 10256 12847 10290
rect 12909 10256 12915 10290
rect 12981 10256 12983 10290
rect 13017 10256 13019 10290
rect 13085 10256 13091 10290
rect 13153 10256 13163 10290
rect 13221 10256 13235 10290
rect 13289 10256 13307 10290
rect 13357 10256 13379 10290
rect 13425 10256 13451 10290
rect 13493 10256 13523 10290
rect 13561 10256 13595 10290
rect 13629 10256 13817 10290
rect 1177 10214 13817 10256
rect 13968 34680 14361 34706
rect 13968 34646 14120 34680
rect 14154 34672 14361 34680
rect 14154 34646 14297 34672
rect 13968 34638 14297 34646
rect 14331 34638 14361 34672
rect 13968 34608 14361 34638
rect 13968 34574 14120 34608
rect 14154 34604 14361 34608
rect 14154 34574 14297 34604
rect 13968 34570 14297 34574
rect 14331 34570 14361 34604
rect 13968 34536 14361 34570
rect 13968 34502 14120 34536
rect 14154 34502 14297 34536
rect 14331 34502 14361 34536
rect 13968 34468 14361 34502
rect 13968 34464 14297 34468
rect 13968 34430 14120 34464
rect 14154 34434 14297 34464
rect 14331 34434 14361 34468
rect 14154 34430 14361 34434
rect 13968 34400 14361 34430
rect 13968 34392 14297 34400
rect 13968 34358 14120 34392
rect 14154 34366 14297 34392
rect 14331 34366 14361 34400
rect 14154 34358 14361 34366
rect 13968 34332 14361 34358
rect 13968 34320 14297 34332
rect 13968 34286 14120 34320
rect 14154 34298 14297 34320
rect 14331 34298 14361 34332
rect 14154 34286 14361 34298
rect 13968 34264 14361 34286
rect 13968 34248 14297 34264
rect 13968 34214 14120 34248
rect 14154 34230 14297 34248
rect 14331 34230 14361 34264
rect 14154 34214 14361 34230
rect 13968 34196 14361 34214
rect 13968 34176 14297 34196
rect 13968 34142 14120 34176
rect 14154 34162 14297 34176
rect 14331 34162 14361 34196
rect 14154 34142 14361 34162
rect 13968 34128 14361 34142
rect 13968 34104 14297 34128
rect 13968 34070 14120 34104
rect 14154 34094 14297 34104
rect 14331 34094 14361 34128
rect 14154 34070 14361 34094
rect 13968 34060 14361 34070
rect 13968 34032 14297 34060
rect 13968 33998 14120 34032
rect 14154 34026 14297 34032
rect 14331 34026 14361 34060
rect 14154 33998 14361 34026
rect 13968 33992 14361 33998
rect 13968 33960 14297 33992
rect 13968 33926 14120 33960
rect 14154 33958 14297 33960
rect 14331 33958 14361 33992
rect 14154 33926 14361 33958
rect 13968 33924 14361 33926
rect 13968 33890 14297 33924
rect 14331 33890 14361 33924
rect 13968 33888 14361 33890
rect 13968 33854 14120 33888
rect 14154 33856 14361 33888
rect 14154 33854 14297 33856
rect 13968 33822 14297 33854
rect 14331 33822 14361 33856
rect 13968 33816 14361 33822
rect 13968 33782 14120 33816
rect 14154 33788 14361 33816
rect 14154 33782 14297 33788
rect 13968 33754 14297 33782
rect 14331 33754 14361 33788
rect 13968 33744 14361 33754
rect 13968 33710 14120 33744
rect 14154 33720 14361 33744
rect 14154 33710 14297 33720
rect 13968 33686 14297 33710
rect 14331 33686 14361 33720
rect 13968 33672 14361 33686
rect 13968 33638 14120 33672
rect 14154 33652 14361 33672
rect 14154 33638 14297 33652
rect 13968 33618 14297 33638
rect 14331 33618 14361 33652
rect 13968 33600 14361 33618
rect 13968 33566 14120 33600
rect 14154 33584 14361 33600
rect 14154 33566 14297 33584
rect 13968 33550 14297 33566
rect 14331 33550 14361 33584
rect 13968 33528 14361 33550
rect 13968 33494 14120 33528
rect 14154 33516 14361 33528
rect 14154 33494 14297 33516
rect 13968 33482 14297 33494
rect 14331 33482 14361 33516
rect 13968 33456 14361 33482
rect 13968 33422 14120 33456
rect 14154 33448 14361 33456
rect 14154 33422 14297 33448
rect 13968 33414 14297 33422
rect 14331 33414 14361 33448
rect 13968 33384 14361 33414
rect 13968 33350 14120 33384
rect 14154 33380 14361 33384
rect 14154 33350 14297 33380
rect 13968 33346 14297 33350
rect 14331 33346 14361 33380
rect 13968 33312 14361 33346
rect 13968 33278 14120 33312
rect 14154 33278 14297 33312
rect 14331 33278 14361 33312
rect 13968 33244 14361 33278
rect 13968 33240 14297 33244
rect 13968 33206 14120 33240
rect 14154 33210 14297 33240
rect 14331 33210 14361 33244
rect 14154 33206 14361 33210
rect 13968 33176 14361 33206
rect 13968 33168 14297 33176
rect 13968 33134 14120 33168
rect 14154 33142 14297 33168
rect 14331 33142 14361 33176
rect 14154 33134 14361 33142
rect 13968 33108 14361 33134
rect 13968 33096 14297 33108
rect 13968 33062 14120 33096
rect 14154 33074 14297 33096
rect 14331 33074 14361 33108
rect 14154 33062 14361 33074
rect 13968 33040 14361 33062
rect 13968 33024 14297 33040
rect 13968 32990 14120 33024
rect 14154 33006 14297 33024
rect 14331 33006 14361 33040
rect 14154 32990 14361 33006
rect 13968 32972 14361 32990
rect 13968 32952 14297 32972
rect 13968 32918 14120 32952
rect 14154 32938 14297 32952
rect 14331 32938 14361 32972
rect 14154 32918 14361 32938
rect 13968 32904 14361 32918
rect 13968 32880 14297 32904
rect 13968 32846 14120 32880
rect 14154 32870 14297 32880
rect 14331 32870 14361 32904
rect 14154 32846 14361 32870
rect 13968 32836 14361 32846
rect 13968 32808 14297 32836
rect 13968 32774 14120 32808
rect 14154 32802 14297 32808
rect 14331 32802 14361 32836
rect 14154 32774 14361 32802
rect 13968 32768 14361 32774
rect 13968 32736 14297 32768
rect 13968 32702 14120 32736
rect 14154 32734 14297 32736
rect 14331 32734 14361 32768
rect 14154 32702 14361 32734
rect 13968 32700 14361 32702
rect 13968 32666 14297 32700
rect 14331 32666 14361 32700
rect 13968 32664 14361 32666
rect 13968 32630 14120 32664
rect 14154 32632 14361 32664
rect 14154 32630 14297 32632
rect 13968 32598 14297 32630
rect 14331 32598 14361 32632
rect 13968 32592 14361 32598
rect 13968 32558 14120 32592
rect 14154 32564 14361 32592
rect 14154 32558 14297 32564
rect 13968 32530 14297 32558
rect 14331 32530 14361 32564
rect 13968 32520 14361 32530
rect 13968 32486 14120 32520
rect 14154 32496 14361 32520
rect 14154 32486 14297 32496
rect 13968 32462 14297 32486
rect 14331 32462 14361 32496
rect 13968 32448 14361 32462
rect 13968 32414 14120 32448
rect 14154 32428 14361 32448
rect 14154 32414 14297 32428
rect 13968 32394 14297 32414
rect 14331 32394 14361 32428
rect 13968 32376 14361 32394
rect 13968 32342 14120 32376
rect 14154 32360 14361 32376
rect 14154 32342 14297 32360
rect 13968 32326 14297 32342
rect 14331 32326 14361 32360
rect 13968 32304 14361 32326
rect 13968 32270 14120 32304
rect 14154 32292 14361 32304
rect 14154 32270 14297 32292
rect 13968 32258 14297 32270
rect 14331 32258 14361 32292
rect 13968 32232 14361 32258
rect 13968 32198 14120 32232
rect 14154 32224 14361 32232
rect 14154 32198 14297 32224
rect 13968 32190 14297 32198
rect 14331 32190 14361 32224
rect 13968 32160 14361 32190
rect 13968 32126 14120 32160
rect 14154 32156 14361 32160
rect 14154 32126 14297 32156
rect 13968 32122 14297 32126
rect 14331 32122 14361 32156
rect 13968 32088 14361 32122
rect 13968 32054 14120 32088
rect 14154 32054 14297 32088
rect 14331 32054 14361 32088
rect 13968 32020 14361 32054
rect 13968 32016 14297 32020
rect 13968 31982 14120 32016
rect 14154 31986 14297 32016
rect 14331 31986 14361 32020
rect 14154 31982 14361 31986
rect 13968 31952 14361 31982
rect 13968 31944 14297 31952
rect 13968 31910 14120 31944
rect 14154 31918 14297 31944
rect 14331 31918 14361 31952
rect 14154 31910 14361 31918
rect 13968 31884 14361 31910
rect 13968 31872 14297 31884
rect 13968 31838 14120 31872
rect 14154 31850 14297 31872
rect 14331 31850 14361 31884
rect 14154 31838 14361 31850
rect 13968 31816 14361 31838
rect 13968 31800 14297 31816
rect 13968 31766 14120 31800
rect 14154 31782 14297 31800
rect 14331 31782 14361 31816
rect 14154 31766 14361 31782
rect 13968 31748 14361 31766
rect 13968 31728 14297 31748
rect 13968 31694 14120 31728
rect 14154 31714 14297 31728
rect 14331 31714 14361 31748
rect 14154 31694 14361 31714
rect 13968 31680 14361 31694
rect 13968 31656 14297 31680
rect 13968 31622 14120 31656
rect 14154 31646 14297 31656
rect 14331 31646 14361 31680
rect 14154 31622 14361 31646
rect 13968 31612 14361 31622
rect 13968 31584 14297 31612
rect 13968 31550 14120 31584
rect 14154 31578 14297 31584
rect 14331 31578 14361 31612
rect 14154 31550 14361 31578
rect 13968 31544 14361 31550
rect 13968 31512 14297 31544
rect 13968 31478 14120 31512
rect 14154 31510 14297 31512
rect 14331 31510 14361 31544
rect 14154 31478 14361 31510
rect 13968 31476 14361 31478
rect 13968 31442 14297 31476
rect 14331 31442 14361 31476
rect 13968 31440 14361 31442
rect 13968 31406 14120 31440
rect 14154 31408 14361 31440
rect 14154 31406 14297 31408
rect 13968 31374 14297 31406
rect 14331 31374 14361 31408
rect 13968 31368 14361 31374
rect 13968 31334 14120 31368
rect 14154 31340 14361 31368
rect 14154 31334 14297 31340
rect 13968 31306 14297 31334
rect 14331 31306 14361 31340
rect 13968 31296 14361 31306
rect 13968 31262 14120 31296
rect 14154 31272 14361 31296
rect 14154 31262 14297 31272
rect 13968 31238 14297 31262
rect 14331 31238 14361 31272
rect 13968 31224 14361 31238
rect 13968 31190 14120 31224
rect 14154 31204 14361 31224
rect 14154 31190 14297 31204
rect 13968 31170 14297 31190
rect 14331 31170 14361 31204
rect 13968 31152 14361 31170
rect 13968 31118 14120 31152
rect 14154 31136 14361 31152
rect 14154 31118 14297 31136
rect 13968 31102 14297 31118
rect 14331 31102 14361 31136
rect 13968 31080 14361 31102
rect 13968 31046 14120 31080
rect 14154 31068 14361 31080
rect 14154 31046 14297 31068
rect 13968 31034 14297 31046
rect 14331 31034 14361 31068
rect 13968 31008 14361 31034
rect 13968 30974 14120 31008
rect 14154 31000 14361 31008
rect 14154 30974 14297 31000
rect 13968 30966 14297 30974
rect 14331 30966 14361 31000
rect 13968 30936 14361 30966
rect 13968 30902 14120 30936
rect 14154 30932 14361 30936
rect 14154 30902 14297 30932
rect 13968 30898 14297 30902
rect 14331 30898 14361 30932
rect 13968 30864 14361 30898
rect 13968 30830 14120 30864
rect 14154 30830 14297 30864
rect 14331 30830 14361 30864
rect 13968 30796 14361 30830
rect 13968 30792 14297 30796
rect 13968 30758 14120 30792
rect 14154 30762 14297 30792
rect 14331 30762 14361 30796
rect 14154 30758 14361 30762
rect 13968 30728 14361 30758
rect 13968 30720 14297 30728
rect 13968 30686 14120 30720
rect 14154 30694 14297 30720
rect 14331 30694 14361 30728
rect 14154 30686 14361 30694
rect 13968 30660 14361 30686
rect 13968 30648 14297 30660
rect 13968 30614 14120 30648
rect 14154 30626 14297 30648
rect 14331 30626 14361 30660
rect 14154 30614 14361 30626
rect 13968 30592 14361 30614
rect 13968 30576 14297 30592
rect 13968 30542 14120 30576
rect 14154 30558 14297 30576
rect 14331 30558 14361 30592
rect 14154 30542 14361 30558
rect 13968 30524 14361 30542
rect 13968 30504 14297 30524
rect 13968 30470 14120 30504
rect 14154 30490 14297 30504
rect 14331 30490 14361 30524
rect 14154 30470 14361 30490
rect 13968 30456 14361 30470
rect 13968 30432 14297 30456
rect 13968 30398 14120 30432
rect 14154 30422 14297 30432
rect 14331 30422 14361 30456
rect 14154 30398 14361 30422
rect 13968 30388 14361 30398
rect 13968 30360 14297 30388
rect 13968 30326 14120 30360
rect 14154 30354 14297 30360
rect 14331 30354 14361 30388
rect 14154 30326 14361 30354
rect 13968 30320 14361 30326
rect 13968 30288 14297 30320
rect 13968 30254 14120 30288
rect 14154 30286 14297 30288
rect 14331 30286 14361 30320
rect 14154 30254 14361 30286
rect 13968 30252 14361 30254
rect 13968 30218 14297 30252
rect 14331 30218 14361 30252
rect 13968 30216 14361 30218
rect 13968 30182 14120 30216
rect 14154 30184 14361 30216
rect 14154 30182 14297 30184
rect 13968 30150 14297 30182
rect 14331 30150 14361 30184
rect 13968 30144 14361 30150
rect 13968 30110 14120 30144
rect 14154 30116 14361 30144
rect 14154 30110 14297 30116
rect 13968 30082 14297 30110
rect 14331 30082 14361 30116
rect 13968 30072 14361 30082
rect 13968 30038 14120 30072
rect 14154 30048 14361 30072
rect 14154 30038 14297 30048
rect 13968 30014 14297 30038
rect 14331 30014 14361 30048
rect 13968 30000 14361 30014
rect 13968 29966 14120 30000
rect 14154 29980 14361 30000
rect 14154 29966 14297 29980
rect 13968 29946 14297 29966
rect 14331 29946 14361 29980
rect 13968 29928 14361 29946
rect 13968 29894 14120 29928
rect 14154 29912 14361 29928
rect 14154 29894 14297 29912
rect 13968 29878 14297 29894
rect 14331 29878 14361 29912
rect 13968 29856 14361 29878
rect 13968 29822 14120 29856
rect 14154 29844 14361 29856
rect 14154 29822 14297 29844
rect 13968 29810 14297 29822
rect 14331 29810 14361 29844
rect 13968 29784 14361 29810
rect 13968 29750 14120 29784
rect 14154 29776 14361 29784
rect 14154 29750 14297 29776
rect 13968 29742 14297 29750
rect 14331 29742 14361 29776
rect 13968 29712 14361 29742
rect 13968 29678 14120 29712
rect 14154 29708 14361 29712
rect 14154 29678 14297 29708
rect 13968 29674 14297 29678
rect 14331 29674 14361 29708
rect 13968 29640 14361 29674
rect 13968 29606 14120 29640
rect 14154 29606 14297 29640
rect 14331 29606 14361 29640
rect 13968 29572 14361 29606
rect 13968 29568 14297 29572
rect 13968 29534 14120 29568
rect 14154 29538 14297 29568
rect 14331 29538 14361 29572
rect 14154 29534 14361 29538
rect 13968 29504 14361 29534
rect 13968 29496 14297 29504
rect 13968 29462 14120 29496
rect 14154 29470 14297 29496
rect 14331 29470 14361 29504
rect 14154 29462 14361 29470
rect 13968 29436 14361 29462
rect 13968 29424 14297 29436
rect 13968 29390 14120 29424
rect 14154 29402 14297 29424
rect 14331 29402 14361 29436
rect 14154 29390 14361 29402
rect 13968 29368 14361 29390
rect 13968 29352 14297 29368
rect 13968 29318 14120 29352
rect 14154 29334 14297 29352
rect 14331 29334 14361 29368
rect 14154 29318 14361 29334
rect 13968 29300 14361 29318
rect 13968 29280 14297 29300
rect 13968 29246 14120 29280
rect 14154 29266 14297 29280
rect 14331 29266 14361 29300
rect 14154 29246 14361 29266
rect 13968 29232 14361 29246
rect 13968 29208 14297 29232
rect 13968 29174 14120 29208
rect 14154 29198 14297 29208
rect 14331 29198 14361 29232
rect 14154 29174 14361 29198
rect 13968 29164 14361 29174
rect 13968 29136 14297 29164
rect 13968 29102 14120 29136
rect 14154 29130 14297 29136
rect 14331 29130 14361 29164
rect 14154 29102 14361 29130
rect 13968 29096 14361 29102
rect 13968 29064 14297 29096
rect 13968 29030 14120 29064
rect 14154 29062 14297 29064
rect 14331 29062 14361 29096
rect 14154 29030 14361 29062
rect 13968 29028 14361 29030
rect 13968 28994 14297 29028
rect 14331 28994 14361 29028
rect 13968 28992 14361 28994
rect 13968 28958 14120 28992
rect 14154 28960 14361 28992
rect 14154 28958 14297 28960
rect 13968 28926 14297 28958
rect 14331 28926 14361 28960
rect 13968 28920 14361 28926
rect 13968 28886 14120 28920
rect 14154 28892 14361 28920
rect 14154 28886 14297 28892
rect 13968 28858 14297 28886
rect 14331 28858 14361 28892
rect 13968 28848 14361 28858
rect 13968 28814 14120 28848
rect 14154 28824 14361 28848
rect 14154 28814 14297 28824
rect 13968 28790 14297 28814
rect 14331 28790 14361 28824
rect 13968 28776 14361 28790
rect 13968 28742 14120 28776
rect 14154 28756 14361 28776
rect 14154 28742 14297 28756
rect 13968 28722 14297 28742
rect 14331 28722 14361 28756
rect 13968 28704 14361 28722
rect 13968 28670 14120 28704
rect 14154 28688 14361 28704
rect 14154 28670 14297 28688
rect 13968 28654 14297 28670
rect 14331 28654 14361 28688
rect 13968 28632 14361 28654
rect 13968 28598 14120 28632
rect 14154 28620 14361 28632
rect 14154 28598 14297 28620
rect 13968 28586 14297 28598
rect 14331 28586 14361 28620
rect 13968 28560 14361 28586
rect 13968 28526 14120 28560
rect 14154 28552 14361 28560
rect 14154 28526 14297 28552
rect 13968 28518 14297 28526
rect 14331 28518 14361 28552
rect 13968 28488 14361 28518
rect 13968 28454 14120 28488
rect 14154 28484 14361 28488
rect 14154 28454 14297 28484
rect 13968 28450 14297 28454
rect 14331 28450 14361 28484
rect 13968 28416 14361 28450
rect 13968 28382 14120 28416
rect 14154 28382 14297 28416
rect 14331 28382 14361 28416
rect 13968 28348 14361 28382
rect 13968 28344 14297 28348
rect 13968 28310 14120 28344
rect 14154 28314 14297 28344
rect 14331 28314 14361 28348
rect 14154 28310 14361 28314
rect 13968 28280 14361 28310
rect 13968 28272 14297 28280
rect 13968 28238 14120 28272
rect 14154 28246 14297 28272
rect 14331 28246 14361 28280
rect 14154 28238 14361 28246
rect 13968 28212 14361 28238
rect 13968 28200 14297 28212
rect 13968 28166 14120 28200
rect 14154 28178 14297 28200
rect 14331 28178 14361 28212
rect 14154 28166 14361 28178
rect 13968 28144 14361 28166
rect 13968 28128 14297 28144
rect 13968 28094 14120 28128
rect 14154 28110 14297 28128
rect 14331 28110 14361 28144
rect 14154 28094 14361 28110
rect 13968 28076 14361 28094
rect 13968 28056 14297 28076
rect 13968 28022 14120 28056
rect 14154 28042 14297 28056
rect 14331 28042 14361 28076
rect 14154 28022 14361 28042
rect 13968 28008 14361 28022
rect 13968 27984 14297 28008
rect 13968 27950 14120 27984
rect 14154 27974 14297 27984
rect 14331 27974 14361 28008
rect 14154 27950 14361 27974
rect 13968 27940 14361 27950
rect 13968 27912 14297 27940
rect 13968 27878 14120 27912
rect 14154 27906 14297 27912
rect 14331 27906 14361 27940
rect 14154 27878 14361 27906
rect 13968 27872 14361 27878
rect 13968 27840 14297 27872
rect 13968 27806 14120 27840
rect 14154 27838 14297 27840
rect 14331 27838 14361 27872
rect 14154 27806 14361 27838
rect 13968 27804 14361 27806
rect 13968 27770 14297 27804
rect 14331 27770 14361 27804
rect 13968 27768 14361 27770
rect 13968 27734 14120 27768
rect 14154 27736 14361 27768
rect 14154 27734 14297 27736
rect 13968 27702 14297 27734
rect 14331 27702 14361 27736
rect 13968 27696 14361 27702
rect 13968 27662 14120 27696
rect 14154 27668 14361 27696
rect 14154 27662 14297 27668
rect 13968 27634 14297 27662
rect 14331 27634 14361 27668
rect 13968 27624 14361 27634
rect 13968 27590 14120 27624
rect 14154 27600 14361 27624
rect 14154 27590 14297 27600
rect 13968 27566 14297 27590
rect 14331 27566 14361 27600
rect 13968 27552 14361 27566
rect 13968 27518 14120 27552
rect 14154 27532 14361 27552
rect 14154 27518 14297 27532
rect 13968 27498 14297 27518
rect 14331 27498 14361 27532
rect 13968 27480 14361 27498
rect 13968 27446 14120 27480
rect 14154 27464 14361 27480
rect 14154 27446 14297 27464
rect 13968 27430 14297 27446
rect 14331 27430 14361 27464
rect 13968 27408 14361 27430
rect 13968 27374 14120 27408
rect 14154 27396 14361 27408
rect 14154 27374 14297 27396
rect 13968 27362 14297 27374
rect 14331 27362 14361 27396
rect 13968 27336 14361 27362
rect 13968 27302 14120 27336
rect 14154 27328 14361 27336
rect 14154 27302 14297 27328
rect 13968 27294 14297 27302
rect 14331 27294 14361 27328
rect 13968 27264 14361 27294
rect 13968 27230 14120 27264
rect 14154 27260 14361 27264
rect 14154 27230 14297 27260
rect 13968 27226 14297 27230
rect 14331 27226 14361 27260
rect 13968 27192 14361 27226
rect 13968 27158 14120 27192
rect 14154 27158 14297 27192
rect 14331 27158 14361 27192
rect 13968 27124 14361 27158
rect 13968 27120 14297 27124
rect 13968 27086 14120 27120
rect 14154 27090 14297 27120
rect 14331 27090 14361 27124
rect 14154 27086 14361 27090
rect 13968 27056 14361 27086
rect 13968 27048 14297 27056
rect 13968 27014 14120 27048
rect 14154 27022 14297 27048
rect 14331 27022 14361 27056
rect 14154 27014 14361 27022
rect 13968 26988 14361 27014
rect 13968 26976 14297 26988
rect 13968 26942 14120 26976
rect 14154 26954 14297 26976
rect 14331 26954 14361 26988
rect 14154 26942 14361 26954
rect 13968 26920 14361 26942
rect 13968 26904 14297 26920
rect 13968 26870 14120 26904
rect 14154 26886 14297 26904
rect 14331 26886 14361 26920
rect 14154 26870 14361 26886
rect 13968 26852 14361 26870
rect 13968 26832 14297 26852
rect 13968 26798 14120 26832
rect 14154 26818 14297 26832
rect 14331 26818 14361 26852
rect 14154 26798 14361 26818
rect 13968 26784 14361 26798
rect 13968 26760 14297 26784
rect 13968 26726 14120 26760
rect 14154 26750 14297 26760
rect 14331 26750 14361 26784
rect 14154 26726 14361 26750
rect 13968 26716 14361 26726
rect 13968 26688 14297 26716
rect 13968 26654 14120 26688
rect 14154 26682 14297 26688
rect 14331 26682 14361 26716
rect 14154 26654 14361 26682
rect 13968 26648 14361 26654
rect 13968 26616 14297 26648
rect 13968 26582 14120 26616
rect 14154 26614 14297 26616
rect 14331 26614 14361 26648
rect 14154 26582 14361 26614
rect 13968 26580 14361 26582
rect 13968 26546 14297 26580
rect 14331 26546 14361 26580
rect 13968 26544 14361 26546
rect 13968 26510 14120 26544
rect 14154 26512 14361 26544
rect 14154 26510 14297 26512
rect 13968 26478 14297 26510
rect 14331 26478 14361 26512
rect 13968 26472 14361 26478
rect 13968 26438 14120 26472
rect 14154 26444 14361 26472
rect 14154 26438 14297 26444
rect 13968 26410 14297 26438
rect 14331 26410 14361 26444
rect 13968 26400 14361 26410
rect 13968 26366 14120 26400
rect 14154 26376 14361 26400
rect 14154 26366 14297 26376
rect 13968 26342 14297 26366
rect 14331 26342 14361 26376
rect 13968 26328 14361 26342
rect 13968 26294 14120 26328
rect 14154 26308 14361 26328
rect 14154 26294 14297 26308
rect 13968 26274 14297 26294
rect 14331 26274 14361 26308
rect 13968 26256 14361 26274
rect 13968 26222 14120 26256
rect 14154 26240 14361 26256
rect 14154 26222 14297 26240
rect 13968 26206 14297 26222
rect 14331 26206 14361 26240
rect 13968 26184 14361 26206
rect 13968 26150 14120 26184
rect 14154 26172 14361 26184
rect 14154 26150 14297 26172
rect 13968 26138 14297 26150
rect 14331 26138 14361 26172
rect 13968 26112 14361 26138
rect 13968 26078 14120 26112
rect 14154 26104 14361 26112
rect 14154 26078 14297 26104
rect 13968 26070 14297 26078
rect 14331 26070 14361 26104
rect 13968 26040 14361 26070
rect 13968 26006 14120 26040
rect 14154 26036 14361 26040
rect 14154 26006 14297 26036
rect 13968 26002 14297 26006
rect 14331 26002 14361 26036
rect 13968 25968 14361 26002
rect 13968 25934 14120 25968
rect 14154 25934 14297 25968
rect 14331 25934 14361 25968
rect 13968 25900 14361 25934
rect 13968 25896 14297 25900
rect 13968 25862 14120 25896
rect 14154 25866 14297 25896
rect 14331 25866 14361 25900
rect 14154 25862 14361 25866
rect 13968 25832 14361 25862
rect 13968 25824 14297 25832
rect 13968 25790 14120 25824
rect 14154 25798 14297 25824
rect 14331 25798 14361 25832
rect 14154 25790 14361 25798
rect 13968 25764 14361 25790
rect 13968 25752 14297 25764
rect 13968 25718 14120 25752
rect 14154 25730 14297 25752
rect 14331 25730 14361 25764
rect 14154 25718 14361 25730
rect 13968 25696 14361 25718
rect 13968 25680 14297 25696
rect 13968 25646 14120 25680
rect 14154 25662 14297 25680
rect 14331 25662 14361 25696
rect 14154 25646 14361 25662
rect 13968 25628 14361 25646
rect 13968 25608 14297 25628
rect 13968 25574 14120 25608
rect 14154 25594 14297 25608
rect 14331 25594 14361 25628
rect 14154 25574 14361 25594
rect 13968 25560 14361 25574
rect 13968 25536 14297 25560
rect 13968 25502 14120 25536
rect 14154 25526 14297 25536
rect 14331 25526 14361 25560
rect 14154 25502 14361 25526
rect 13968 25492 14361 25502
rect 13968 25464 14297 25492
rect 13968 25430 14120 25464
rect 14154 25458 14297 25464
rect 14331 25458 14361 25492
rect 14154 25430 14361 25458
rect 13968 25424 14361 25430
rect 13968 25392 14297 25424
rect 13968 25358 14120 25392
rect 14154 25390 14297 25392
rect 14331 25390 14361 25424
rect 14154 25358 14361 25390
rect 13968 25356 14361 25358
rect 13968 25322 14297 25356
rect 14331 25322 14361 25356
rect 13968 25320 14361 25322
rect 13968 25286 14120 25320
rect 14154 25288 14361 25320
rect 14154 25286 14297 25288
rect 13968 25254 14297 25286
rect 14331 25254 14361 25288
rect 13968 25248 14361 25254
rect 13968 25214 14120 25248
rect 14154 25220 14361 25248
rect 14154 25214 14297 25220
rect 13968 25186 14297 25214
rect 14331 25186 14361 25220
rect 13968 25176 14361 25186
rect 13968 25142 14120 25176
rect 14154 25152 14361 25176
rect 14154 25142 14297 25152
rect 13968 25118 14297 25142
rect 14331 25118 14361 25152
rect 13968 25104 14361 25118
rect 13968 25070 14120 25104
rect 14154 25084 14361 25104
rect 14154 25070 14297 25084
rect 13968 25050 14297 25070
rect 14331 25050 14361 25084
rect 13968 25032 14361 25050
rect 13968 24998 14120 25032
rect 14154 25016 14361 25032
rect 14154 24998 14297 25016
rect 13968 24982 14297 24998
rect 14331 24982 14361 25016
rect 13968 24960 14361 24982
rect 13968 24926 14120 24960
rect 14154 24948 14361 24960
rect 14154 24926 14297 24948
rect 13968 24914 14297 24926
rect 14331 24914 14361 24948
rect 13968 24888 14361 24914
rect 13968 24854 14120 24888
rect 14154 24880 14361 24888
rect 14154 24854 14297 24880
rect 13968 24846 14297 24854
rect 14331 24846 14361 24880
rect 13968 24816 14361 24846
rect 13968 24782 14120 24816
rect 14154 24812 14361 24816
rect 14154 24782 14297 24812
rect 13968 24778 14297 24782
rect 14331 24778 14361 24812
rect 13968 24744 14361 24778
rect 13968 24710 14120 24744
rect 14154 24710 14297 24744
rect 14331 24710 14361 24744
rect 13968 24676 14361 24710
rect 13968 24672 14297 24676
rect 13968 24638 14120 24672
rect 14154 24642 14297 24672
rect 14331 24642 14361 24676
rect 14154 24638 14361 24642
rect 13968 24608 14361 24638
rect 13968 24600 14297 24608
rect 13968 24566 14120 24600
rect 14154 24574 14297 24600
rect 14331 24574 14361 24608
rect 14154 24566 14361 24574
rect 13968 24540 14361 24566
rect 13968 24528 14297 24540
rect 13968 24494 14120 24528
rect 14154 24506 14297 24528
rect 14331 24506 14361 24540
rect 14154 24494 14361 24506
rect 13968 24472 14361 24494
rect 13968 24456 14297 24472
rect 13968 24422 14120 24456
rect 14154 24438 14297 24456
rect 14331 24438 14361 24472
rect 14154 24422 14361 24438
rect 13968 24404 14361 24422
rect 13968 24384 14297 24404
rect 13968 24350 14120 24384
rect 14154 24370 14297 24384
rect 14331 24370 14361 24404
rect 14154 24350 14361 24370
rect 13968 24336 14361 24350
rect 13968 24312 14297 24336
rect 13968 24278 14120 24312
rect 14154 24302 14297 24312
rect 14331 24302 14361 24336
rect 14154 24278 14361 24302
rect 13968 24268 14361 24278
rect 13968 24240 14297 24268
rect 13968 24206 14120 24240
rect 14154 24234 14297 24240
rect 14331 24234 14361 24268
rect 14154 24206 14361 24234
rect 13968 24200 14361 24206
rect 13968 24168 14297 24200
rect 13968 24134 14120 24168
rect 14154 24166 14297 24168
rect 14331 24166 14361 24200
rect 14154 24134 14361 24166
rect 13968 24132 14361 24134
rect 13968 24098 14297 24132
rect 14331 24098 14361 24132
rect 13968 24096 14361 24098
rect 13968 24062 14120 24096
rect 14154 24064 14361 24096
rect 14154 24062 14297 24064
rect 13968 24030 14297 24062
rect 14331 24030 14361 24064
rect 13968 24024 14361 24030
rect 13968 23990 14120 24024
rect 14154 23996 14361 24024
rect 14154 23990 14297 23996
rect 13968 23962 14297 23990
rect 14331 23962 14361 23996
rect 13968 23952 14361 23962
rect 13968 23918 14120 23952
rect 14154 23928 14361 23952
rect 14154 23918 14297 23928
rect 13968 23894 14297 23918
rect 14331 23894 14361 23928
rect 13968 23880 14361 23894
rect 13968 23846 14120 23880
rect 14154 23860 14361 23880
rect 14154 23846 14297 23860
rect 13968 23826 14297 23846
rect 14331 23826 14361 23860
rect 13968 23808 14361 23826
rect 13968 23774 14120 23808
rect 14154 23792 14361 23808
rect 14154 23774 14297 23792
rect 13968 23758 14297 23774
rect 14331 23758 14361 23792
rect 13968 23736 14361 23758
rect 13968 23702 14120 23736
rect 14154 23724 14361 23736
rect 14154 23702 14297 23724
rect 13968 23690 14297 23702
rect 14331 23690 14361 23724
rect 13968 23664 14361 23690
rect 13968 23630 14120 23664
rect 14154 23656 14361 23664
rect 14154 23630 14297 23656
rect 13968 23622 14297 23630
rect 14331 23622 14361 23656
rect 13968 23592 14361 23622
rect 13968 23558 14120 23592
rect 14154 23588 14361 23592
rect 14154 23558 14297 23588
rect 13968 23554 14297 23558
rect 14331 23554 14361 23588
rect 13968 23520 14361 23554
rect 13968 23486 14120 23520
rect 14154 23486 14297 23520
rect 14331 23486 14361 23520
rect 13968 23452 14361 23486
rect 13968 23448 14297 23452
rect 13968 23414 14120 23448
rect 14154 23418 14297 23448
rect 14331 23418 14361 23452
rect 14154 23414 14361 23418
rect 13968 23384 14361 23414
rect 13968 23376 14297 23384
rect 13968 23342 14120 23376
rect 14154 23350 14297 23376
rect 14331 23350 14361 23384
rect 14154 23342 14361 23350
rect 13968 23316 14361 23342
rect 13968 23304 14297 23316
rect 13968 23270 14120 23304
rect 14154 23282 14297 23304
rect 14331 23282 14361 23316
rect 14154 23270 14361 23282
rect 13968 23248 14361 23270
rect 13968 23232 14297 23248
rect 13968 23198 14120 23232
rect 14154 23214 14297 23232
rect 14331 23214 14361 23248
rect 14154 23198 14361 23214
rect 13968 23180 14361 23198
rect 13968 23160 14297 23180
rect 13968 23126 14120 23160
rect 14154 23146 14297 23160
rect 14331 23146 14361 23180
rect 14154 23126 14361 23146
rect 13968 23112 14361 23126
rect 13968 23088 14297 23112
rect 13968 23054 14120 23088
rect 14154 23078 14297 23088
rect 14331 23078 14361 23112
rect 14154 23054 14361 23078
rect 13968 23044 14361 23054
rect 13968 23016 14297 23044
rect 13968 22982 14120 23016
rect 14154 23010 14297 23016
rect 14331 23010 14361 23044
rect 14154 22982 14361 23010
rect 13968 22976 14361 22982
rect 13968 22944 14297 22976
rect 13968 22910 14120 22944
rect 14154 22942 14297 22944
rect 14331 22942 14361 22976
rect 14154 22910 14361 22942
rect 13968 22908 14361 22910
rect 13968 22874 14297 22908
rect 14331 22874 14361 22908
rect 13968 22872 14361 22874
rect 13968 22838 14120 22872
rect 14154 22840 14361 22872
rect 14154 22838 14297 22840
rect 13968 22806 14297 22838
rect 14331 22806 14361 22840
rect 13968 22800 14361 22806
rect 13968 22766 14120 22800
rect 14154 22772 14361 22800
rect 14154 22766 14297 22772
rect 13968 22738 14297 22766
rect 14331 22738 14361 22772
rect 13968 22728 14361 22738
rect 13968 22694 14120 22728
rect 14154 22704 14361 22728
rect 14154 22694 14297 22704
rect 13968 22670 14297 22694
rect 14331 22670 14361 22704
rect 13968 22656 14361 22670
rect 13968 22622 14120 22656
rect 14154 22636 14361 22656
rect 14154 22622 14297 22636
rect 13968 22602 14297 22622
rect 14331 22602 14361 22636
rect 13968 22584 14361 22602
rect 13968 22550 14120 22584
rect 14154 22568 14361 22584
rect 14154 22550 14297 22568
rect 13968 22534 14297 22550
rect 14331 22534 14361 22568
rect 13968 22512 14361 22534
rect 13968 22478 14120 22512
rect 14154 22500 14361 22512
rect 14154 22478 14297 22500
rect 13968 22466 14297 22478
rect 14331 22466 14361 22500
rect 13968 22440 14361 22466
rect 13968 22406 14120 22440
rect 14154 22432 14361 22440
rect 14154 22406 14297 22432
rect 13968 22398 14297 22406
rect 14331 22398 14361 22432
rect 13968 22368 14361 22398
rect 13968 22334 14120 22368
rect 14154 22364 14361 22368
rect 14154 22334 14297 22364
rect 13968 22330 14297 22334
rect 14331 22330 14361 22364
rect 13968 22296 14361 22330
rect 13968 22262 14120 22296
rect 14154 22262 14297 22296
rect 14331 22262 14361 22296
rect 13968 22228 14361 22262
rect 13968 22224 14297 22228
rect 13968 22190 14120 22224
rect 14154 22194 14297 22224
rect 14331 22194 14361 22228
rect 14154 22190 14361 22194
rect 13968 22160 14361 22190
rect 13968 22152 14297 22160
rect 13968 22118 14120 22152
rect 14154 22126 14297 22152
rect 14331 22126 14361 22160
rect 14154 22118 14361 22126
rect 13968 22092 14361 22118
rect 13968 22080 14297 22092
rect 13968 22046 14120 22080
rect 14154 22058 14297 22080
rect 14331 22058 14361 22092
rect 14154 22046 14361 22058
rect 13968 22024 14361 22046
rect 13968 22008 14297 22024
rect 13968 21974 14120 22008
rect 14154 21990 14297 22008
rect 14331 21990 14361 22024
rect 14154 21974 14361 21990
rect 13968 21956 14361 21974
rect 13968 21936 14297 21956
rect 13968 21902 14120 21936
rect 14154 21922 14297 21936
rect 14331 21922 14361 21956
rect 14154 21902 14361 21922
rect 13968 21888 14361 21902
rect 13968 21864 14297 21888
rect 13968 21830 14120 21864
rect 14154 21854 14297 21864
rect 14331 21854 14361 21888
rect 14154 21830 14361 21854
rect 13968 21820 14361 21830
rect 13968 21792 14297 21820
rect 13968 21758 14120 21792
rect 14154 21786 14297 21792
rect 14331 21786 14361 21820
rect 14154 21758 14361 21786
rect 13968 21752 14361 21758
rect 13968 21720 14297 21752
rect 13968 21686 14120 21720
rect 14154 21718 14297 21720
rect 14331 21718 14361 21752
rect 14154 21686 14361 21718
rect 13968 21684 14361 21686
rect 13968 21650 14297 21684
rect 14331 21650 14361 21684
rect 13968 21648 14361 21650
rect 13968 21614 14120 21648
rect 14154 21616 14361 21648
rect 14154 21614 14297 21616
rect 13968 21582 14297 21614
rect 14331 21582 14361 21616
rect 13968 21576 14361 21582
rect 13968 21542 14120 21576
rect 14154 21548 14361 21576
rect 14154 21542 14297 21548
rect 13968 21514 14297 21542
rect 14331 21514 14361 21548
rect 13968 21504 14361 21514
rect 13968 21470 14120 21504
rect 14154 21480 14361 21504
rect 14154 21470 14297 21480
rect 13968 21446 14297 21470
rect 14331 21446 14361 21480
rect 13968 21432 14361 21446
rect 13968 21398 14120 21432
rect 14154 21412 14361 21432
rect 14154 21398 14297 21412
rect 13968 21378 14297 21398
rect 14331 21378 14361 21412
rect 13968 21360 14361 21378
rect 13968 21326 14120 21360
rect 14154 21344 14361 21360
rect 14154 21326 14297 21344
rect 13968 21310 14297 21326
rect 14331 21310 14361 21344
rect 13968 21288 14361 21310
rect 13968 21254 14120 21288
rect 14154 21276 14361 21288
rect 14154 21254 14297 21276
rect 13968 21242 14297 21254
rect 14331 21242 14361 21276
rect 13968 21216 14361 21242
rect 13968 21182 14120 21216
rect 14154 21208 14361 21216
rect 14154 21182 14297 21208
rect 13968 21174 14297 21182
rect 14331 21174 14361 21208
rect 13968 21144 14361 21174
rect 13968 21110 14120 21144
rect 14154 21140 14361 21144
rect 14154 21110 14297 21140
rect 13968 21106 14297 21110
rect 14331 21106 14361 21140
rect 13968 21072 14361 21106
rect 13968 21038 14120 21072
rect 14154 21038 14297 21072
rect 14331 21038 14361 21072
rect 13968 21004 14361 21038
rect 13968 21000 14297 21004
rect 13968 20966 14120 21000
rect 14154 20970 14297 21000
rect 14331 20970 14361 21004
rect 14154 20966 14361 20970
rect 13968 20936 14361 20966
rect 13968 20928 14297 20936
rect 13968 20894 14120 20928
rect 14154 20902 14297 20928
rect 14331 20902 14361 20936
rect 14154 20894 14361 20902
rect 13968 20868 14361 20894
rect 13968 20856 14297 20868
rect 13968 20822 14120 20856
rect 14154 20834 14297 20856
rect 14331 20834 14361 20868
rect 14154 20822 14361 20834
rect 13968 20800 14361 20822
rect 13968 20784 14297 20800
rect 13968 20750 14120 20784
rect 14154 20766 14297 20784
rect 14331 20766 14361 20800
rect 14154 20750 14361 20766
rect 13968 20732 14361 20750
rect 13968 20712 14297 20732
rect 13968 20678 14120 20712
rect 14154 20698 14297 20712
rect 14331 20698 14361 20732
rect 14154 20678 14361 20698
rect 13968 20664 14361 20678
rect 13968 20640 14297 20664
rect 13968 20606 14120 20640
rect 14154 20630 14297 20640
rect 14331 20630 14361 20664
rect 14154 20606 14361 20630
rect 13968 20596 14361 20606
rect 13968 20568 14297 20596
rect 13968 20534 14120 20568
rect 14154 20562 14297 20568
rect 14331 20562 14361 20596
rect 14154 20534 14361 20562
rect 13968 20528 14361 20534
rect 13968 20496 14297 20528
rect 13968 20462 14120 20496
rect 14154 20494 14297 20496
rect 14331 20494 14361 20528
rect 14154 20462 14361 20494
rect 13968 20460 14361 20462
rect 13968 20426 14297 20460
rect 14331 20426 14361 20460
rect 13968 20424 14361 20426
rect 13968 20390 14120 20424
rect 14154 20392 14361 20424
rect 14154 20390 14297 20392
rect 13968 20358 14297 20390
rect 14331 20358 14361 20392
rect 13968 20352 14361 20358
rect 13968 20318 14120 20352
rect 14154 20324 14361 20352
rect 14154 20318 14297 20324
rect 13968 20290 14297 20318
rect 14331 20290 14361 20324
rect 13968 20280 14361 20290
rect 13968 20246 14120 20280
rect 14154 20256 14361 20280
rect 14154 20246 14297 20256
rect 13968 20222 14297 20246
rect 14331 20222 14361 20256
rect 13968 20208 14361 20222
rect 13968 20174 14120 20208
rect 14154 20188 14361 20208
rect 14154 20174 14297 20188
rect 13968 20154 14297 20174
rect 14331 20154 14361 20188
rect 13968 20136 14361 20154
rect 13968 20102 14120 20136
rect 14154 20120 14361 20136
rect 14154 20102 14297 20120
rect 13968 20086 14297 20102
rect 14331 20086 14361 20120
rect 13968 20064 14361 20086
rect 13968 20030 14120 20064
rect 14154 20052 14361 20064
rect 14154 20030 14297 20052
rect 13968 20018 14297 20030
rect 14331 20018 14361 20052
rect 13968 19992 14361 20018
rect 13968 19958 14120 19992
rect 14154 19984 14361 19992
rect 14154 19958 14297 19984
rect 13968 19950 14297 19958
rect 14331 19950 14361 19984
rect 13968 19920 14361 19950
rect 13968 19886 14120 19920
rect 14154 19916 14361 19920
rect 14154 19886 14297 19916
rect 13968 19882 14297 19886
rect 14331 19882 14361 19916
rect 13968 19848 14361 19882
rect 13968 19814 14120 19848
rect 14154 19814 14297 19848
rect 14331 19814 14361 19848
rect 13968 19780 14361 19814
rect 13968 19776 14297 19780
rect 13968 19742 14120 19776
rect 14154 19746 14297 19776
rect 14331 19746 14361 19780
rect 14154 19742 14361 19746
rect 13968 19712 14361 19742
rect 13968 19704 14297 19712
rect 13968 19670 14120 19704
rect 14154 19678 14297 19704
rect 14331 19678 14361 19712
rect 14154 19670 14361 19678
rect 13968 19644 14361 19670
rect 13968 19632 14297 19644
rect 13968 19598 14120 19632
rect 14154 19610 14297 19632
rect 14331 19610 14361 19644
rect 14154 19598 14361 19610
rect 13968 19576 14361 19598
rect 13968 19560 14297 19576
rect 13968 19526 14120 19560
rect 14154 19542 14297 19560
rect 14331 19542 14361 19576
rect 14154 19526 14361 19542
rect 13968 19508 14361 19526
rect 13968 19488 14297 19508
rect 13968 19454 14120 19488
rect 14154 19474 14297 19488
rect 14331 19474 14361 19508
rect 14154 19454 14361 19474
rect 13968 19440 14361 19454
rect 13968 19416 14297 19440
rect 13968 19382 14120 19416
rect 14154 19406 14297 19416
rect 14331 19406 14361 19440
rect 14154 19382 14361 19406
rect 13968 19372 14361 19382
rect 13968 19344 14297 19372
rect 13968 19310 14120 19344
rect 14154 19338 14297 19344
rect 14331 19338 14361 19372
rect 14154 19310 14361 19338
rect 13968 19304 14361 19310
rect 13968 19272 14297 19304
rect 13968 19238 14120 19272
rect 14154 19270 14297 19272
rect 14331 19270 14361 19304
rect 14154 19238 14361 19270
rect 13968 19236 14361 19238
rect 13968 19202 14297 19236
rect 14331 19202 14361 19236
rect 13968 19200 14361 19202
rect 13968 19166 14120 19200
rect 14154 19168 14361 19200
rect 14154 19166 14297 19168
rect 13968 19134 14297 19166
rect 14331 19134 14361 19168
rect 13968 19128 14361 19134
rect 13968 19094 14120 19128
rect 14154 19100 14361 19128
rect 14154 19094 14297 19100
rect 13968 19066 14297 19094
rect 14331 19066 14361 19100
rect 13968 19056 14361 19066
rect 13968 19022 14120 19056
rect 14154 19032 14361 19056
rect 14154 19022 14297 19032
rect 13968 18998 14297 19022
rect 14331 18998 14361 19032
rect 13968 18984 14361 18998
rect 13968 18950 14120 18984
rect 14154 18964 14361 18984
rect 14154 18950 14297 18964
rect 13968 18930 14297 18950
rect 14331 18930 14361 18964
rect 13968 18912 14361 18930
rect 13968 18878 14120 18912
rect 14154 18896 14361 18912
rect 14154 18878 14297 18896
rect 13968 18862 14297 18878
rect 14331 18862 14361 18896
rect 13968 18840 14361 18862
rect 13968 18806 14120 18840
rect 14154 18828 14361 18840
rect 14154 18806 14297 18828
rect 13968 18794 14297 18806
rect 14331 18794 14361 18828
rect 13968 18768 14361 18794
rect 13968 18734 14120 18768
rect 14154 18760 14361 18768
rect 14154 18734 14297 18760
rect 13968 18726 14297 18734
rect 14331 18726 14361 18760
rect 13968 18696 14361 18726
rect 13968 18662 14120 18696
rect 14154 18692 14361 18696
rect 14154 18662 14297 18692
rect 13968 18658 14297 18662
rect 14331 18658 14361 18692
rect 13968 18624 14361 18658
rect 13968 18590 14120 18624
rect 14154 18590 14297 18624
rect 14331 18590 14361 18624
rect 13968 18556 14361 18590
rect 13968 18552 14297 18556
rect 13968 18518 14120 18552
rect 14154 18522 14297 18552
rect 14331 18522 14361 18556
rect 14154 18518 14361 18522
rect 13968 18488 14361 18518
rect 13968 18480 14297 18488
rect 13968 18446 14120 18480
rect 14154 18454 14297 18480
rect 14331 18454 14361 18488
rect 14154 18446 14361 18454
rect 13968 18420 14361 18446
rect 13968 18408 14297 18420
rect 13968 18374 14120 18408
rect 14154 18386 14297 18408
rect 14331 18386 14361 18420
rect 14154 18374 14361 18386
rect 13968 18352 14361 18374
rect 13968 18336 14297 18352
rect 13968 18302 14120 18336
rect 14154 18318 14297 18336
rect 14331 18318 14361 18352
rect 14154 18302 14361 18318
rect 13968 18284 14361 18302
rect 13968 18264 14297 18284
rect 13968 18230 14120 18264
rect 14154 18250 14297 18264
rect 14331 18250 14361 18284
rect 14154 18230 14361 18250
rect 13968 18216 14361 18230
rect 13968 18192 14297 18216
rect 13968 18158 14120 18192
rect 14154 18182 14297 18192
rect 14331 18182 14361 18216
rect 14154 18158 14361 18182
rect 13968 18148 14361 18158
rect 13968 18120 14297 18148
rect 13968 18086 14120 18120
rect 14154 18114 14297 18120
rect 14331 18114 14361 18148
rect 14154 18086 14361 18114
rect 13968 18080 14361 18086
rect 13968 18048 14297 18080
rect 13968 18014 14120 18048
rect 14154 18046 14297 18048
rect 14331 18046 14361 18080
rect 14154 18014 14361 18046
rect 13968 18012 14361 18014
rect 13968 17978 14297 18012
rect 14331 17978 14361 18012
rect 13968 17976 14361 17978
rect 13968 17942 14120 17976
rect 14154 17944 14361 17976
rect 14154 17942 14297 17944
rect 13968 17910 14297 17942
rect 14331 17910 14361 17944
rect 13968 17904 14361 17910
rect 13968 17870 14120 17904
rect 14154 17876 14361 17904
rect 14154 17870 14297 17876
rect 13968 17842 14297 17870
rect 14331 17842 14361 17876
rect 13968 17832 14361 17842
rect 13968 17798 14120 17832
rect 14154 17808 14361 17832
rect 14154 17798 14297 17808
rect 13968 17774 14297 17798
rect 14331 17774 14361 17808
rect 13968 17760 14361 17774
rect 13968 17726 14120 17760
rect 14154 17740 14361 17760
rect 14154 17726 14297 17740
rect 13968 17706 14297 17726
rect 14331 17706 14361 17740
rect 13968 17688 14361 17706
rect 13968 17654 14120 17688
rect 14154 17672 14361 17688
rect 14154 17654 14297 17672
rect 13968 17638 14297 17654
rect 14331 17638 14361 17672
rect 13968 17616 14361 17638
rect 13968 17582 14120 17616
rect 14154 17604 14361 17616
rect 14154 17582 14297 17604
rect 13968 17570 14297 17582
rect 14331 17570 14361 17604
rect 13968 17544 14361 17570
rect 13968 17510 14120 17544
rect 14154 17536 14361 17544
rect 14154 17510 14297 17536
rect 13968 17502 14297 17510
rect 14331 17502 14361 17536
rect 13968 17472 14361 17502
rect 13968 17438 14120 17472
rect 14154 17468 14361 17472
rect 14154 17438 14297 17468
rect 13968 17434 14297 17438
rect 14331 17434 14361 17468
rect 13968 17400 14361 17434
rect 13968 17366 14120 17400
rect 14154 17366 14297 17400
rect 14331 17366 14361 17400
rect 13968 17332 14361 17366
rect 13968 17328 14297 17332
rect 13968 17294 14120 17328
rect 14154 17298 14297 17328
rect 14331 17298 14361 17332
rect 14154 17294 14361 17298
rect 13968 17264 14361 17294
rect 13968 17256 14297 17264
rect 13968 17222 14120 17256
rect 14154 17230 14297 17256
rect 14331 17230 14361 17264
rect 14154 17222 14361 17230
rect 13968 17196 14361 17222
rect 13968 17184 14297 17196
rect 13968 17150 14120 17184
rect 14154 17162 14297 17184
rect 14331 17162 14361 17196
rect 14154 17150 14361 17162
rect 13968 17128 14361 17150
rect 13968 17112 14297 17128
rect 13968 17078 14120 17112
rect 14154 17094 14297 17112
rect 14331 17094 14361 17128
rect 14154 17078 14361 17094
rect 13968 17060 14361 17078
rect 13968 17040 14297 17060
rect 13968 17006 14120 17040
rect 14154 17026 14297 17040
rect 14331 17026 14361 17060
rect 14154 17006 14361 17026
rect 13968 16992 14361 17006
rect 13968 16968 14297 16992
rect 13968 16934 14120 16968
rect 14154 16958 14297 16968
rect 14331 16958 14361 16992
rect 14154 16934 14361 16958
rect 13968 16924 14361 16934
rect 13968 16896 14297 16924
rect 13968 16862 14120 16896
rect 14154 16890 14297 16896
rect 14331 16890 14361 16924
rect 14154 16862 14361 16890
rect 13968 16856 14361 16862
rect 13968 16824 14297 16856
rect 13968 16790 14120 16824
rect 14154 16822 14297 16824
rect 14331 16822 14361 16856
rect 14154 16790 14361 16822
rect 13968 16788 14361 16790
rect 13968 16754 14297 16788
rect 14331 16754 14361 16788
rect 13968 16752 14361 16754
rect 13968 16718 14120 16752
rect 14154 16720 14361 16752
rect 14154 16718 14297 16720
rect 13968 16686 14297 16718
rect 14331 16686 14361 16720
rect 13968 16680 14361 16686
rect 13968 16646 14120 16680
rect 14154 16652 14361 16680
rect 14154 16646 14297 16652
rect 13968 16618 14297 16646
rect 14331 16618 14361 16652
rect 13968 16608 14361 16618
rect 13968 16574 14120 16608
rect 14154 16584 14361 16608
rect 14154 16574 14297 16584
rect 13968 16550 14297 16574
rect 14331 16550 14361 16584
rect 13968 16536 14361 16550
rect 13968 16502 14120 16536
rect 14154 16516 14361 16536
rect 14154 16502 14297 16516
rect 13968 16482 14297 16502
rect 14331 16482 14361 16516
rect 13968 16464 14361 16482
rect 13968 16430 14120 16464
rect 14154 16448 14361 16464
rect 14154 16430 14297 16448
rect 13968 16414 14297 16430
rect 14331 16414 14361 16448
rect 13968 16392 14361 16414
rect 13968 16358 14120 16392
rect 14154 16380 14361 16392
rect 14154 16358 14297 16380
rect 13968 16346 14297 16358
rect 14331 16346 14361 16380
rect 13968 16320 14361 16346
rect 13968 16286 14120 16320
rect 14154 16312 14361 16320
rect 14154 16286 14297 16312
rect 13968 16278 14297 16286
rect 14331 16278 14361 16312
rect 13968 16248 14361 16278
rect 13968 16214 14120 16248
rect 14154 16244 14361 16248
rect 14154 16214 14297 16244
rect 13968 16210 14297 16214
rect 14331 16210 14361 16244
rect 13968 16176 14361 16210
rect 13968 16142 14120 16176
rect 14154 16142 14297 16176
rect 14331 16142 14361 16176
rect 13968 16108 14361 16142
rect 13968 16104 14297 16108
rect 13968 16070 14120 16104
rect 14154 16074 14297 16104
rect 14331 16074 14361 16108
rect 14154 16070 14361 16074
rect 13968 16040 14361 16070
rect 13968 16032 14297 16040
rect 13968 15998 14120 16032
rect 14154 16006 14297 16032
rect 14331 16006 14361 16040
rect 14154 15998 14361 16006
rect 13968 15972 14361 15998
rect 13968 15960 14297 15972
rect 13968 15926 14120 15960
rect 14154 15938 14297 15960
rect 14331 15938 14361 15972
rect 14154 15926 14361 15938
rect 13968 15904 14361 15926
rect 13968 15888 14297 15904
rect 13968 15854 14120 15888
rect 14154 15870 14297 15888
rect 14331 15870 14361 15904
rect 14154 15854 14361 15870
rect 13968 15836 14361 15854
rect 13968 15816 14297 15836
rect 13968 15782 14120 15816
rect 14154 15802 14297 15816
rect 14331 15802 14361 15836
rect 14154 15782 14361 15802
rect 13968 15768 14361 15782
rect 13968 15744 14297 15768
rect 13968 15710 14120 15744
rect 14154 15734 14297 15744
rect 14331 15734 14361 15768
rect 14154 15710 14361 15734
rect 13968 15700 14361 15710
rect 13968 15672 14297 15700
rect 13968 15638 14120 15672
rect 14154 15666 14297 15672
rect 14331 15666 14361 15700
rect 14154 15638 14361 15666
rect 13968 15632 14361 15638
rect 13968 15600 14297 15632
rect 13968 15566 14120 15600
rect 14154 15598 14297 15600
rect 14331 15598 14361 15632
rect 14154 15566 14361 15598
rect 13968 15564 14361 15566
rect 13968 15530 14297 15564
rect 14331 15530 14361 15564
rect 13968 15528 14361 15530
rect 13968 15494 14120 15528
rect 14154 15496 14361 15528
rect 14154 15494 14297 15496
rect 13968 15462 14297 15494
rect 14331 15462 14361 15496
rect 13968 15456 14361 15462
rect 13968 15422 14120 15456
rect 14154 15428 14361 15456
rect 14154 15422 14297 15428
rect 13968 15394 14297 15422
rect 14331 15394 14361 15428
rect 13968 15384 14361 15394
rect 13968 15350 14120 15384
rect 14154 15360 14361 15384
rect 14154 15350 14297 15360
rect 13968 15326 14297 15350
rect 14331 15326 14361 15360
rect 13968 15312 14361 15326
rect 13968 15278 14120 15312
rect 14154 15292 14361 15312
rect 14154 15278 14297 15292
rect 13968 15258 14297 15278
rect 14331 15258 14361 15292
rect 13968 15240 14361 15258
rect 13968 15206 14120 15240
rect 14154 15224 14361 15240
rect 14154 15206 14297 15224
rect 13968 15190 14297 15206
rect 14331 15190 14361 15224
rect 13968 15168 14361 15190
rect 13968 15134 14120 15168
rect 14154 15156 14361 15168
rect 14154 15134 14297 15156
rect 13968 15122 14297 15134
rect 14331 15122 14361 15156
rect 13968 15096 14361 15122
rect 13968 15062 14120 15096
rect 14154 15088 14361 15096
rect 14154 15062 14297 15088
rect 13968 15054 14297 15062
rect 14331 15054 14361 15088
rect 13968 15024 14361 15054
rect 13968 14990 14120 15024
rect 14154 15020 14361 15024
rect 14154 14990 14297 15020
rect 13968 14986 14297 14990
rect 14331 14986 14361 15020
rect 13968 14952 14361 14986
rect 13968 14918 14120 14952
rect 14154 14918 14297 14952
rect 14331 14918 14361 14952
rect 13968 14884 14361 14918
rect 13968 14880 14297 14884
rect 13968 14846 14120 14880
rect 14154 14850 14297 14880
rect 14331 14850 14361 14884
rect 14154 14846 14361 14850
rect 13968 14816 14361 14846
rect 13968 14808 14297 14816
rect 13968 14774 14120 14808
rect 14154 14782 14297 14808
rect 14331 14782 14361 14816
rect 14154 14774 14361 14782
rect 13968 14748 14361 14774
rect 13968 14736 14297 14748
rect 13968 14702 14120 14736
rect 14154 14714 14297 14736
rect 14331 14714 14361 14748
rect 14154 14702 14361 14714
rect 13968 14680 14361 14702
rect 13968 14664 14297 14680
rect 13968 14630 14120 14664
rect 14154 14646 14297 14664
rect 14331 14646 14361 14680
rect 14154 14630 14361 14646
rect 13968 14612 14361 14630
rect 13968 14592 14297 14612
rect 13968 14558 14120 14592
rect 14154 14578 14297 14592
rect 14331 14578 14361 14612
rect 14154 14558 14361 14578
rect 13968 14544 14361 14558
rect 13968 14520 14297 14544
rect 13968 14486 14120 14520
rect 14154 14510 14297 14520
rect 14331 14510 14361 14544
rect 14154 14486 14361 14510
rect 13968 14476 14361 14486
rect 13968 14448 14297 14476
rect 13968 14414 14120 14448
rect 14154 14442 14297 14448
rect 14331 14442 14361 14476
rect 14154 14414 14361 14442
rect 13968 14408 14361 14414
rect 13968 14376 14297 14408
rect 13968 14342 14120 14376
rect 14154 14374 14297 14376
rect 14331 14374 14361 14408
rect 14154 14342 14361 14374
rect 13968 14340 14361 14342
rect 13968 14306 14297 14340
rect 14331 14306 14361 14340
rect 13968 14304 14361 14306
rect 13968 14270 14120 14304
rect 14154 14272 14361 14304
rect 14154 14270 14297 14272
rect 13968 14238 14297 14270
rect 14331 14238 14361 14272
rect 13968 14232 14361 14238
rect 13968 14198 14120 14232
rect 14154 14204 14361 14232
rect 14154 14198 14297 14204
rect 13968 14170 14297 14198
rect 14331 14170 14361 14204
rect 13968 14160 14361 14170
rect 13968 14126 14120 14160
rect 14154 14136 14361 14160
rect 14154 14126 14297 14136
rect 13968 14102 14297 14126
rect 14331 14102 14361 14136
rect 13968 14088 14361 14102
rect 13968 14054 14120 14088
rect 14154 14068 14361 14088
rect 14154 14054 14297 14068
rect 13968 14034 14297 14054
rect 14331 14034 14361 14068
rect 13968 14016 14361 14034
rect 13968 13982 14120 14016
rect 14154 14000 14361 14016
rect 14154 13982 14297 14000
rect 13968 13966 14297 13982
rect 14331 13966 14361 14000
rect 13968 13944 14361 13966
rect 13968 13910 14120 13944
rect 14154 13932 14361 13944
rect 14154 13910 14297 13932
rect 13968 13898 14297 13910
rect 14331 13898 14361 13932
rect 13968 13872 14361 13898
rect 13968 13838 14120 13872
rect 14154 13864 14361 13872
rect 14154 13838 14297 13864
rect 13968 13830 14297 13838
rect 14331 13830 14361 13864
rect 13968 13800 14361 13830
rect 13968 13766 14120 13800
rect 14154 13796 14361 13800
rect 14154 13766 14297 13796
rect 13968 13762 14297 13766
rect 14331 13762 14361 13796
rect 13968 13728 14361 13762
rect 13968 13694 14120 13728
rect 14154 13694 14297 13728
rect 14331 13694 14361 13728
rect 13968 13660 14361 13694
rect 13968 13656 14297 13660
rect 13968 13622 14120 13656
rect 14154 13626 14297 13656
rect 14331 13626 14361 13660
rect 14154 13622 14361 13626
rect 13968 13592 14361 13622
rect 13968 13584 14297 13592
rect 13968 13550 14120 13584
rect 14154 13558 14297 13584
rect 14331 13558 14361 13592
rect 14154 13550 14361 13558
rect 13968 13524 14361 13550
rect 13968 13512 14297 13524
rect 13968 13478 14120 13512
rect 14154 13490 14297 13512
rect 14331 13490 14361 13524
rect 14154 13478 14361 13490
rect 13968 13456 14361 13478
rect 13968 13440 14297 13456
rect 13968 13406 14120 13440
rect 14154 13422 14297 13440
rect 14331 13422 14361 13456
rect 14154 13406 14361 13422
rect 13968 13388 14361 13406
rect 13968 13368 14297 13388
rect 13968 13334 14120 13368
rect 14154 13354 14297 13368
rect 14331 13354 14361 13388
rect 14154 13334 14361 13354
rect 13968 13320 14361 13334
rect 13968 13296 14297 13320
rect 13968 13262 14120 13296
rect 14154 13286 14297 13296
rect 14331 13286 14361 13320
rect 14154 13262 14361 13286
rect 13968 13252 14361 13262
rect 13968 13224 14297 13252
rect 13968 13190 14120 13224
rect 14154 13218 14297 13224
rect 14331 13218 14361 13252
rect 14154 13190 14361 13218
rect 13968 13184 14361 13190
rect 13968 13152 14297 13184
rect 13968 13118 14120 13152
rect 14154 13150 14297 13152
rect 14331 13150 14361 13184
rect 14154 13118 14361 13150
rect 13968 13116 14361 13118
rect 13968 13082 14297 13116
rect 14331 13082 14361 13116
rect 13968 13080 14361 13082
rect 13968 13046 14120 13080
rect 14154 13048 14361 13080
rect 14154 13046 14297 13048
rect 13968 13014 14297 13046
rect 14331 13014 14361 13048
rect 13968 13008 14361 13014
rect 13968 12974 14120 13008
rect 14154 12980 14361 13008
rect 14154 12974 14297 12980
rect 13968 12946 14297 12974
rect 14331 12946 14361 12980
rect 13968 12936 14361 12946
rect 13968 12902 14120 12936
rect 14154 12912 14361 12936
rect 14154 12902 14297 12912
rect 13968 12878 14297 12902
rect 14331 12878 14361 12912
rect 13968 12864 14361 12878
rect 13968 12830 14120 12864
rect 14154 12844 14361 12864
rect 14154 12830 14297 12844
rect 13968 12810 14297 12830
rect 14331 12810 14361 12844
rect 13968 12792 14361 12810
rect 13968 12758 14120 12792
rect 14154 12776 14361 12792
rect 14154 12758 14297 12776
rect 13968 12742 14297 12758
rect 14331 12742 14361 12776
rect 13968 12720 14361 12742
rect 13968 12686 14120 12720
rect 14154 12708 14361 12720
rect 14154 12686 14297 12708
rect 13968 12674 14297 12686
rect 14331 12674 14361 12708
rect 13968 12648 14361 12674
rect 13968 12614 14120 12648
rect 14154 12640 14361 12648
rect 14154 12614 14297 12640
rect 13968 12606 14297 12614
rect 14331 12606 14361 12640
rect 13968 12576 14361 12606
rect 13968 12542 14120 12576
rect 14154 12572 14361 12576
rect 14154 12542 14297 12572
rect 13968 12538 14297 12542
rect 14331 12538 14361 12572
rect 13968 12504 14361 12538
rect 13968 12470 14120 12504
rect 14154 12470 14297 12504
rect 14331 12470 14361 12504
rect 13968 12436 14361 12470
rect 13968 12432 14297 12436
rect 13968 12398 14120 12432
rect 14154 12402 14297 12432
rect 14331 12402 14361 12436
rect 14154 12398 14361 12402
rect 13968 12368 14361 12398
rect 13968 12360 14297 12368
rect 13968 12326 14120 12360
rect 14154 12334 14297 12360
rect 14331 12334 14361 12368
rect 14154 12326 14361 12334
rect 13968 12300 14361 12326
rect 13968 12288 14297 12300
rect 13968 12254 14120 12288
rect 14154 12266 14297 12288
rect 14331 12266 14361 12300
rect 14154 12254 14361 12266
rect 13968 12232 14361 12254
rect 13968 12216 14297 12232
rect 13968 12182 14120 12216
rect 14154 12198 14297 12216
rect 14331 12198 14361 12232
rect 14154 12182 14361 12198
rect 13968 12164 14361 12182
rect 13968 12144 14297 12164
rect 13968 12110 14120 12144
rect 14154 12130 14297 12144
rect 14331 12130 14361 12164
rect 14154 12110 14361 12130
rect 13968 12096 14361 12110
rect 13968 12072 14297 12096
rect 13968 12038 14120 12072
rect 14154 12062 14297 12072
rect 14331 12062 14361 12096
rect 14154 12038 14361 12062
rect 13968 12028 14361 12038
rect 13968 12000 14297 12028
rect 13968 11966 14120 12000
rect 14154 11994 14297 12000
rect 14331 11994 14361 12028
rect 14154 11966 14361 11994
rect 13968 11960 14361 11966
rect 13968 11928 14297 11960
rect 13968 11894 14120 11928
rect 14154 11926 14297 11928
rect 14331 11926 14361 11960
rect 14154 11894 14361 11926
rect 13968 11892 14361 11894
rect 13968 11858 14297 11892
rect 14331 11858 14361 11892
rect 13968 11856 14361 11858
rect 13968 11822 14120 11856
rect 14154 11824 14361 11856
rect 14154 11822 14297 11824
rect 13968 11790 14297 11822
rect 14331 11790 14361 11824
rect 13968 11784 14361 11790
rect 13968 11750 14120 11784
rect 14154 11756 14361 11784
rect 14154 11750 14297 11756
rect 13968 11722 14297 11750
rect 14331 11722 14361 11756
rect 13968 11712 14361 11722
rect 13968 11678 14120 11712
rect 14154 11688 14361 11712
rect 14154 11678 14297 11688
rect 13968 11654 14297 11678
rect 14331 11654 14361 11688
rect 13968 11640 14361 11654
rect 13968 11606 14120 11640
rect 14154 11620 14361 11640
rect 14154 11606 14297 11620
rect 13968 11586 14297 11606
rect 14331 11586 14361 11620
rect 13968 11568 14361 11586
rect 13968 11534 14120 11568
rect 14154 11552 14361 11568
rect 14154 11534 14297 11552
rect 13968 11518 14297 11534
rect 14331 11518 14361 11552
rect 13968 11496 14361 11518
rect 13968 11462 14120 11496
rect 14154 11484 14361 11496
rect 14154 11462 14297 11484
rect 13968 11450 14297 11462
rect 14331 11450 14361 11484
rect 13968 11424 14361 11450
rect 13968 11390 14120 11424
rect 14154 11416 14361 11424
rect 14154 11390 14297 11416
rect 13968 11382 14297 11390
rect 14331 11382 14361 11416
rect 13968 11352 14361 11382
rect 13968 11318 14120 11352
rect 14154 11348 14361 11352
rect 14154 11318 14297 11348
rect 13968 11314 14297 11318
rect 14331 11314 14361 11348
rect 13968 11280 14361 11314
rect 13968 11246 14120 11280
rect 14154 11246 14297 11280
rect 14331 11246 14361 11280
rect 13968 11212 14361 11246
rect 13968 11208 14297 11212
rect 13968 11174 14120 11208
rect 14154 11178 14297 11208
rect 14331 11178 14361 11212
rect 14154 11174 14361 11178
rect 13968 11144 14361 11174
rect 13968 11136 14297 11144
rect 13968 11102 14120 11136
rect 14154 11110 14297 11136
rect 14331 11110 14361 11144
rect 14154 11102 14361 11110
rect 13968 11076 14361 11102
rect 13968 11064 14297 11076
rect 13968 11030 14120 11064
rect 14154 11042 14297 11064
rect 14331 11042 14361 11076
rect 14154 11030 14361 11042
rect 13968 11008 14361 11030
rect 13968 10992 14297 11008
rect 13968 10958 14120 10992
rect 14154 10974 14297 10992
rect 14331 10974 14361 11008
rect 14154 10958 14361 10974
rect 13968 10940 14361 10958
rect 13968 10920 14297 10940
rect 13968 10886 14120 10920
rect 14154 10906 14297 10920
rect 14331 10906 14361 10940
rect 14154 10886 14361 10906
rect 13968 10872 14361 10886
rect 13968 10848 14297 10872
rect 13968 10814 14120 10848
rect 14154 10838 14297 10848
rect 14331 10838 14361 10872
rect 14154 10814 14361 10838
rect 13968 10804 14361 10814
rect 13968 10776 14297 10804
rect 13968 10742 14120 10776
rect 14154 10770 14297 10776
rect 14331 10770 14361 10804
rect 14154 10742 14361 10770
rect 13968 10736 14361 10742
rect 13968 10704 14297 10736
rect 13968 10670 14120 10704
rect 14154 10702 14297 10704
rect 14331 10702 14361 10736
rect 14154 10670 14361 10702
rect 13968 10668 14361 10670
rect 13968 10634 14297 10668
rect 14331 10634 14361 10668
rect 13968 10632 14361 10634
rect 13968 10598 14120 10632
rect 14154 10600 14361 10632
rect 14154 10598 14297 10600
rect 13968 10566 14297 10598
rect 14331 10566 14361 10600
rect 13968 10560 14361 10566
rect 13968 10526 14120 10560
rect 14154 10532 14361 10560
rect 14154 10526 14297 10532
rect 13968 10498 14297 10526
rect 14331 10498 14361 10532
rect 13968 10488 14361 10498
rect 13968 10454 14120 10488
rect 14154 10464 14361 10488
rect 14154 10454 14297 10464
rect 13968 10430 14297 10454
rect 14331 10430 14361 10464
rect 13968 10416 14361 10430
rect 13968 10382 14120 10416
rect 14154 10396 14361 10416
rect 14154 10382 14297 10396
rect 13968 10362 14297 10382
rect 14331 10362 14361 10396
rect 13968 10344 14361 10362
rect 13968 10310 14120 10344
rect 14154 10328 14361 10344
rect 14154 10310 14297 10328
rect 13968 10294 14297 10310
rect 14331 10294 14361 10328
rect 13968 10272 14361 10294
rect 13968 10238 14120 10272
rect 14154 10260 14361 10272
rect 14154 10238 14297 10260
rect 13968 10226 14297 10238
rect 14331 10226 14361 10260
rect 617 10192 814 10207
rect 617 10158 646 10192
rect 680 10173 814 10192
rect 848 10173 1026 10207
rect 680 10158 1026 10173
rect 617 10135 1026 10158
rect 617 10124 814 10135
rect 617 10090 646 10124
rect 680 10101 814 10124
rect 848 10101 1026 10135
rect 680 10093 1026 10101
rect 13968 10200 14361 10226
rect 13968 10166 14120 10200
rect 14154 10192 14361 10200
rect 14154 10166 14297 10192
rect 13968 10158 14297 10166
rect 14331 10158 14361 10192
rect 13968 10128 14361 10158
rect 13968 10094 14120 10128
rect 14154 10124 14361 10128
rect 14154 10094 14297 10124
rect 13968 10093 14297 10094
rect 680 10090 14297 10093
rect 14331 10090 14361 10124
rect 617 10056 14361 10090
rect 617 10022 646 10056
rect 680 10022 14297 10056
rect 14331 10022 14361 10056
rect 617 9988 14361 10022
rect 617 9954 646 9988
rect 680 9954 14297 9988
rect 14331 9954 14361 9988
rect 617 9942 14361 9954
rect 617 9920 912 9942
rect 617 9886 646 9920
rect 680 9908 912 9920
rect 946 9908 984 9942
rect 1018 9908 1056 9942
rect 1090 9908 1128 9942
rect 1162 9908 1200 9942
rect 1234 9908 1272 9942
rect 1306 9908 1344 9942
rect 1378 9908 1416 9942
rect 1450 9908 1488 9942
rect 1522 9908 1560 9942
rect 1594 9908 1632 9942
rect 1666 9908 1704 9942
rect 1738 9908 1776 9942
rect 1810 9908 1848 9942
rect 1882 9908 1920 9942
rect 1954 9908 1992 9942
rect 2026 9908 2064 9942
rect 2098 9908 2136 9942
rect 2170 9908 2208 9942
rect 2242 9908 2280 9942
rect 2314 9908 2352 9942
rect 2386 9908 2424 9942
rect 2458 9908 2496 9942
rect 2530 9908 2568 9942
rect 2602 9908 2640 9942
rect 2674 9908 2712 9942
rect 2746 9908 2784 9942
rect 2818 9908 2856 9942
rect 2890 9908 2928 9942
rect 2962 9908 3000 9942
rect 3034 9908 3072 9942
rect 3106 9908 3144 9942
rect 3178 9908 3216 9942
rect 3250 9908 3288 9942
rect 3322 9908 3360 9942
rect 3394 9908 3432 9942
rect 3466 9908 3504 9942
rect 3538 9908 3576 9942
rect 3610 9908 3648 9942
rect 3682 9908 3720 9942
rect 3754 9908 3792 9942
rect 3826 9908 3864 9942
rect 3898 9908 3936 9942
rect 3970 9908 4008 9942
rect 4042 9908 4080 9942
rect 4114 9908 4152 9942
rect 4186 9908 4224 9942
rect 4258 9908 4296 9942
rect 4330 9908 4368 9942
rect 4402 9908 4440 9942
rect 4474 9908 4512 9942
rect 4546 9908 4584 9942
rect 4618 9908 4656 9942
rect 4690 9908 4728 9942
rect 4762 9908 4800 9942
rect 4834 9908 4872 9942
rect 4906 9908 4944 9942
rect 4978 9908 5016 9942
rect 5050 9908 5088 9942
rect 5122 9908 5160 9942
rect 5194 9908 5232 9942
rect 5266 9908 5304 9942
rect 5338 9908 5376 9942
rect 5410 9908 5448 9942
rect 5482 9908 5520 9942
rect 5554 9908 5592 9942
rect 5626 9908 5664 9942
rect 5698 9908 5736 9942
rect 5770 9908 5808 9942
rect 5842 9908 5880 9942
rect 5914 9908 5952 9942
rect 5986 9908 6024 9942
rect 6058 9908 6096 9942
rect 6130 9908 6168 9942
rect 6202 9908 6240 9942
rect 6274 9908 6312 9942
rect 6346 9908 6384 9942
rect 6418 9908 6456 9942
rect 6490 9908 6528 9942
rect 6562 9908 6600 9942
rect 6634 9908 6672 9942
rect 6706 9908 6744 9942
rect 6778 9908 6816 9942
rect 6850 9908 6888 9942
rect 6922 9908 6960 9942
rect 6994 9908 7032 9942
rect 7066 9908 7104 9942
rect 7138 9908 7176 9942
rect 7210 9908 7248 9942
rect 7282 9908 7320 9942
rect 7354 9908 7392 9942
rect 7426 9908 7464 9942
rect 7498 9908 7536 9942
rect 7570 9908 7608 9942
rect 7642 9908 7680 9942
rect 7714 9908 7752 9942
rect 7786 9908 7824 9942
rect 7858 9908 7896 9942
rect 7930 9908 7968 9942
rect 8002 9908 8040 9942
rect 8074 9908 8112 9942
rect 8146 9908 8184 9942
rect 8218 9908 8256 9942
rect 8290 9908 8328 9942
rect 8362 9908 8400 9942
rect 8434 9908 8472 9942
rect 8506 9908 8544 9942
rect 8578 9908 8616 9942
rect 8650 9908 8688 9942
rect 8722 9908 8760 9942
rect 8794 9908 8832 9942
rect 8866 9908 8904 9942
rect 8938 9908 8976 9942
rect 9010 9908 9048 9942
rect 9082 9908 9120 9942
rect 9154 9908 9192 9942
rect 9226 9908 9264 9942
rect 9298 9908 9336 9942
rect 9370 9908 9408 9942
rect 9442 9908 9480 9942
rect 9514 9908 9552 9942
rect 9586 9908 9624 9942
rect 9658 9908 9696 9942
rect 9730 9908 9768 9942
rect 9802 9908 9840 9942
rect 9874 9908 9912 9942
rect 9946 9908 9984 9942
rect 10018 9908 10056 9942
rect 10090 9908 10128 9942
rect 10162 9908 10200 9942
rect 10234 9908 10272 9942
rect 10306 9908 10344 9942
rect 10378 9908 10416 9942
rect 10450 9908 10488 9942
rect 10522 9908 10560 9942
rect 10594 9908 10632 9942
rect 10666 9908 10704 9942
rect 10738 9908 10776 9942
rect 10810 9908 10848 9942
rect 10882 9908 10920 9942
rect 10954 9908 10992 9942
rect 11026 9908 11064 9942
rect 11098 9908 11136 9942
rect 11170 9908 11208 9942
rect 11242 9908 11280 9942
rect 11314 9908 11352 9942
rect 11386 9908 11424 9942
rect 11458 9908 11496 9942
rect 11530 9908 11568 9942
rect 11602 9908 11640 9942
rect 11674 9908 11712 9942
rect 11746 9908 11784 9942
rect 11818 9908 11856 9942
rect 11890 9908 11928 9942
rect 11962 9908 12000 9942
rect 12034 9908 12072 9942
rect 12106 9908 12144 9942
rect 12178 9908 12216 9942
rect 12250 9908 12288 9942
rect 12322 9908 12360 9942
rect 12394 9908 12432 9942
rect 12466 9908 12504 9942
rect 12538 9908 12576 9942
rect 12610 9908 12648 9942
rect 12682 9908 12720 9942
rect 12754 9908 12792 9942
rect 12826 9908 12864 9942
rect 12898 9908 12936 9942
rect 12970 9908 13008 9942
rect 13042 9908 13080 9942
rect 13114 9908 13152 9942
rect 13186 9908 13224 9942
rect 13258 9908 13296 9942
rect 13330 9908 13368 9942
rect 13402 9908 13440 9942
rect 13474 9908 13512 9942
rect 13546 9908 13584 9942
rect 13618 9908 13656 9942
rect 13690 9908 13728 9942
rect 13762 9908 13800 9942
rect 13834 9908 13872 9942
rect 13906 9908 13944 9942
rect 13978 9908 14016 9942
rect 14050 9920 14361 9942
rect 14050 9908 14297 9920
rect 680 9886 14297 9908
rect 14331 9886 14361 9920
rect 617 9775 14361 9886
rect 617 9741 773 9775
rect 807 9741 841 9775
rect 875 9774 909 9775
rect 943 9774 977 9775
rect 1011 9774 1045 9775
rect 1079 9774 1113 9775
rect 1147 9774 1181 9775
rect 1215 9774 1249 9775
rect 1283 9774 1317 9775
rect 875 9741 883 9774
rect 943 9741 955 9774
rect 1011 9741 1027 9774
rect 1079 9741 1099 9774
rect 1147 9741 1171 9774
rect 1215 9741 1243 9774
rect 1283 9741 1315 9774
rect 1351 9741 1385 9775
rect 1419 9774 1453 9775
rect 1487 9774 1521 9775
rect 1555 9774 1589 9775
rect 1623 9774 1657 9775
rect 1691 9774 1725 9775
rect 1759 9774 1793 9775
rect 1827 9774 1861 9775
rect 1895 9774 1929 9775
rect 1421 9741 1453 9774
rect 1493 9741 1521 9774
rect 1565 9741 1589 9774
rect 1637 9741 1657 9774
rect 1709 9741 1725 9774
rect 1781 9741 1793 9774
rect 1853 9741 1861 9774
rect 1925 9741 1929 9774
rect 1963 9774 1997 9775
rect 617 9740 883 9741
rect 917 9740 955 9741
rect 989 9740 1027 9741
rect 1061 9740 1099 9741
rect 1133 9740 1171 9741
rect 1205 9740 1243 9741
rect 1277 9740 1315 9741
rect 1349 9740 1387 9741
rect 1421 9740 1459 9741
rect 1493 9740 1531 9741
rect 1565 9740 1603 9741
rect 1637 9740 1675 9741
rect 1709 9740 1747 9741
rect 1781 9740 1819 9741
rect 1853 9740 1891 9741
rect 1925 9740 1963 9741
rect 2031 9774 2065 9775
rect 2031 9741 2035 9774
rect 2099 9741 2133 9775
rect 2167 9741 2201 9775
rect 2235 9741 2269 9775
rect 2303 9741 2337 9775
rect 2371 9741 2405 9775
rect 2439 9741 2473 9775
rect 2507 9741 2541 9775
rect 2575 9741 2609 9775
rect 2643 9741 2677 9775
rect 2711 9741 2745 9775
rect 2779 9741 2813 9775
rect 2847 9741 2881 9775
rect 2915 9741 2949 9775
rect 2983 9741 3017 9775
rect 3051 9741 3085 9775
rect 3119 9741 3153 9775
rect 3187 9741 3221 9775
rect 3255 9741 3289 9775
rect 3323 9741 3357 9775
rect 3391 9741 3425 9775
rect 3459 9741 3493 9775
rect 3527 9741 3561 9775
rect 3595 9741 3629 9775
rect 3663 9741 3697 9775
rect 3731 9741 3765 9775
rect 3799 9741 3833 9775
rect 3867 9741 3901 9775
rect 3935 9741 3969 9775
rect 4003 9741 4037 9775
rect 4071 9741 4105 9775
rect 4139 9741 4173 9775
rect 4207 9741 4241 9775
rect 4275 9741 4309 9775
rect 4343 9741 4377 9775
rect 4411 9741 4445 9775
rect 4479 9741 4513 9775
rect 4547 9741 4581 9775
rect 4615 9741 4649 9775
rect 4683 9741 4717 9775
rect 4751 9741 4785 9775
rect 4819 9741 4853 9775
rect 4887 9741 4921 9775
rect 4955 9741 4989 9775
rect 5023 9741 5057 9775
rect 5091 9741 5125 9775
rect 5159 9741 5193 9775
rect 5227 9741 5261 9775
rect 5295 9741 5329 9775
rect 5363 9741 5397 9775
rect 5431 9741 5465 9775
rect 5499 9741 5533 9775
rect 5567 9741 5601 9775
rect 5635 9741 5669 9775
rect 5703 9741 5737 9775
rect 5771 9741 5805 9775
rect 5839 9741 5873 9775
rect 5907 9741 5941 9775
rect 5975 9741 6009 9775
rect 6043 9741 6077 9775
rect 6111 9741 6145 9775
rect 6179 9741 6213 9775
rect 6247 9741 6281 9775
rect 6315 9741 6349 9775
rect 6383 9741 6417 9775
rect 6451 9741 6485 9775
rect 6519 9741 6553 9775
rect 6587 9741 6621 9775
rect 6655 9741 6689 9775
rect 6723 9741 6757 9775
rect 6791 9741 6825 9775
rect 6859 9741 6893 9775
rect 6927 9741 6961 9775
rect 6995 9741 7029 9775
rect 7063 9741 7097 9775
rect 7131 9741 7165 9775
rect 7199 9741 7233 9775
rect 7267 9741 7301 9775
rect 7335 9741 7369 9775
rect 7403 9741 7437 9775
rect 7471 9741 7505 9775
rect 7539 9741 7573 9775
rect 7607 9741 7641 9775
rect 7675 9741 7709 9775
rect 7743 9741 7777 9775
rect 7811 9741 7845 9775
rect 7879 9741 7913 9775
rect 7947 9741 7981 9775
rect 8015 9741 8049 9775
rect 8083 9741 8117 9775
rect 8151 9741 8185 9775
rect 8219 9741 8253 9775
rect 8287 9741 8321 9775
rect 8355 9741 8389 9775
rect 8423 9741 8457 9775
rect 8491 9741 8525 9775
rect 8559 9741 8593 9775
rect 8627 9741 8661 9775
rect 8695 9741 8729 9775
rect 8763 9741 8797 9775
rect 8831 9741 8865 9775
rect 8899 9741 8933 9775
rect 8967 9741 9001 9775
rect 9035 9741 9069 9775
rect 9103 9741 9137 9775
rect 9171 9741 9205 9775
rect 9239 9741 9273 9775
rect 9307 9741 9341 9775
rect 9375 9741 9409 9775
rect 9443 9741 9477 9775
rect 9511 9741 9545 9775
rect 9579 9741 9613 9775
rect 9647 9741 9681 9775
rect 9715 9741 9749 9775
rect 9783 9741 9817 9775
rect 9851 9741 9885 9775
rect 9919 9741 9953 9775
rect 9987 9741 10021 9775
rect 10055 9741 10089 9775
rect 10123 9741 10157 9775
rect 10191 9741 10225 9775
rect 10259 9741 10293 9775
rect 10327 9741 10361 9775
rect 10395 9741 10429 9775
rect 10463 9741 10497 9775
rect 10531 9741 10565 9775
rect 10599 9741 10633 9775
rect 10667 9741 10701 9775
rect 10735 9741 10769 9775
rect 10803 9741 10837 9775
rect 10871 9741 10905 9775
rect 10939 9741 10973 9775
rect 11007 9741 11041 9775
rect 11075 9741 11109 9775
rect 11143 9741 11177 9775
rect 11211 9741 11245 9775
rect 11279 9741 11313 9775
rect 11347 9741 11381 9775
rect 11415 9741 11449 9775
rect 11483 9741 11517 9775
rect 11551 9741 11585 9775
rect 11619 9741 11653 9775
rect 11687 9741 11721 9775
rect 11755 9741 11789 9775
rect 11823 9741 11857 9775
rect 11891 9741 11925 9775
rect 11959 9741 11993 9775
rect 12027 9741 12061 9775
rect 12095 9741 12129 9775
rect 12163 9741 12197 9775
rect 12231 9741 12265 9775
rect 12299 9741 12333 9775
rect 12367 9741 12401 9775
rect 12435 9741 12469 9775
rect 12503 9741 12537 9775
rect 12571 9741 12605 9775
rect 12639 9741 12673 9775
rect 12707 9741 12741 9775
rect 12775 9741 12809 9775
rect 12843 9741 12877 9775
rect 12911 9774 12945 9775
rect 12979 9774 13013 9775
rect 13047 9774 13081 9775
rect 13115 9774 13149 9775
rect 13183 9774 13217 9775
rect 13251 9774 13285 9775
rect 13319 9774 13353 9775
rect 12917 9741 12945 9774
rect 12989 9741 13013 9774
rect 13061 9741 13081 9774
rect 13133 9741 13149 9774
rect 13205 9741 13217 9774
rect 13277 9741 13285 9774
rect 13349 9741 13353 9774
rect 13387 9774 13421 9775
rect 1997 9740 2035 9741
rect 2069 9740 12883 9741
rect 12917 9740 12955 9741
rect 12989 9740 13027 9741
rect 13061 9740 13099 9741
rect 13133 9740 13171 9741
rect 13205 9740 13243 9741
rect 13277 9740 13315 9741
rect 13349 9740 13387 9741
rect 13455 9774 13489 9775
rect 13523 9774 13557 9775
rect 13591 9774 13625 9775
rect 13659 9774 13693 9775
rect 13727 9774 13761 9775
rect 13795 9774 13829 9775
rect 13863 9774 13897 9775
rect 13931 9774 13965 9775
rect 13455 9741 13459 9774
rect 13523 9741 13531 9774
rect 13591 9741 13603 9774
rect 13659 9741 13675 9774
rect 13727 9741 13747 9774
rect 13795 9741 13819 9774
rect 13863 9741 13891 9774
rect 13931 9741 13963 9774
rect 13999 9741 14033 9775
rect 14067 9774 14101 9775
rect 14069 9741 14101 9774
rect 14135 9741 14169 9775
rect 14203 9741 14361 9775
rect 13421 9740 13459 9741
rect 13493 9740 13531 9741
rect 13565 9740 13603 9741
rect 13637 9740 13675 9741
rect 13709 9740 13747 9741
rect 13781 9740 13819 9741
rect 13853 9740 13891 9741
rect 13925 9740 13963 9741
rect 13997 9740 14035 9741
rect 14069 9740 14361 9741
rect 617 9711 14361 9740
rect 14539 36191 14724 36225
rect 14539 36157 14609 36191
rect 14643 36190 14724 36191
rect 14539 36156 14614 36157
rect 14648 36156 14724 36190
rect 14539 36123 14724 36156
rect 14539 36089 14609 36123
rect 14643 36118 14724 36123
rect 14539 36084 14614 36089
rect 14648 36084 14724 36118
rect 14539 36055 14724 36084
rect 14539 36021 14609 36055
rect 14643 36046 14724 36055
rect 14539 36012 14614 36021
rect 14648 36012 14724 36046
rect 14539 35987 14724 36012
rect 14539 35953 14609 35987
rect 14643 35974 14724 35987
rect 14539 35940 14614 35953
rect 14648 35940 14724 35974
rect 14539 35919 14724 35940
rect 14539 35885 14609 35919
rect 14643 35902 14724 35919
rect 14539 35868 14614 35885
rect 14648 35868 14724 35902
rect 14539 35851 14724 35868
rect 14539 35817 14609 35851
rect 14643 35830 14724 35851
rect 14539 35796 14614 35817
rect 14648 35796 14724 35830
rect 14539 35783 14724 35796
rect 14539 35749 14609 35783
rect 14643 35758 14724 35783
rect 14539 35724 14614 35749
rect 14648 35724 14724 35758
rect 14539 35715 14724 35724
rect 14539 35681 14609 35715
rect 14643 35686 14724 35715
rect 14539 35652 14614 35681
rect 14648 35652 14724 35686
rect 14539 35647 14724 35652
rect 14539 35613 14609 35647
rect 14643 35614 14724 35647
rect 14539 35580 14614 35613
rect 14648 35580 14724 35614
rect 14539 35579 14724 35580
rect 14539 35545 14609 35579
rect 14643 35545 14724 35579
rect 14539 35542 14724 35545
rect 14539 35511 14614 35542
rect 14539 35477 14609 35511
rect 14648 35508 14724 35542
rect 14643 35477 14724 35508
rect 14539 35470 14724 35477
rect 14539 35443 14614 35470
rect 14539 35409 14609 35443
rect 14648 35436 14724 35470
rect 14643 35409 14724 35436
rect 14539 35398 14724 35409
rect 14539 35375 14614 35398
rect 14539 35341 14609 35375
rect 14648 35364 14724 35398
rect 14643 35341 14724 35364
rect 14539 35326 14724 35341
rect 14539 35307 14614 35326
rect 14539 35273 14609 35307
rect 14648 35292 14724 35326
rect 14643 35273 14724 35292
rect 14539 35254 14724 35273
rect 14539 35239 14614 35254
rect 14539 35205 14609 35239
rect 14648 35220 14724 35254
rect 14643 35205 14724 35220
rect 14539 35182 14724 35205
rect 14539 35171 14614 35182
rect 14539 35137 14609 35171
rect 14648 35148 14724 35182
rect 14643 35137 14724 35148
rect 14539 35110 14724 35137
rect 14539 35103 14614 35110
rect 14539 35069 14609 35103
rect 14648 35076 14724 35110
rect 14643 35069 14724 35076
rect 14539 35038 14724 35069
rect 14539 35035 14614 35038
rect 14539 35001 14609 35035
rect 14648 35004 14724 35038
rect 14643 35001 14724 35004
rect 14539 34967 14724 35001
rect 14539 34933 14609 34967
rect 14643 34966 14724 34967
rect 14539 34932 14614 34933
rect 14648 34932 14724 34966
rect 14539 34899 14724 34932
rect 14539 34865 14609 34899
rect 14643 34894 14724 34899
rect 14539 34860 14614 34865
rect 14648 34860 14724 34894
rect 14539 34831 14724 34860
rect 14539 34797 14609 34831
rect 14643 34822 14724 34831
rect 14539 34788 14614 34797
rect 14648 34788 14724 34822
rect 14539 34763 14724 34788
rect 14539 34729 14609 34763
rect 14643 34750 14724 34763
rect 14539 34716 14614 34729
rect 14648 34716 14724 34750
rect 14539 34695 14724 34716
rect 14539 34661 14609 34695
rect 14643 34678 14724 34695
rect 14539 34644 14614 34661
rect 14648 34644 14724 34678
rect 14539 34627 14724 34644
rect 14539 34593 14609 34627
rect 14643 34606 14724 34627
rect 14539 34572 14614 34593
rect 14648 34572 14724 34606
rect 14539 34559 14724 34572
rect 14539 34525 14609 34559
rect 14643 34534 14724 34559
rect 14539 34500 14614 34525
rect 14648 34500 14724 34534
rect 14539 34491 14724 34500
rect 14539 34457 14609 34491
rect 14643 34462 14724 34491
rect 14539 34428 14614 34457
rect 14648 34428 14724 34462
rect 14539 34423 14724 34428
rect 14539 34389 14609 34423
rect 14643 34390 14724 34423
rect 14539 34356 14614 34389
rect 14648 34356 14724 34390
rect 14539 34355 14724 34356
rect 14539 34321 14609 34355
rect 14643 34321 14724 34355
rect 14539 34318 14724 34321
rect 14539 34287 14614 34318
rect 14539 34253 14609 34287
rect 14648 34284 14724 34318
rect 14643 34253 14724 34284
rect 14539 34246 14724 34253
rect 14539 34219 14614 34246
rect 14539 34185 14609 34219
rect 14648 34212 14724 34246
rect 14643 34185 14724 34212
rect 14539 34174 14724 34185
rect 14539 34151 14614 34174
rect 14539 34117 14609 34151
rect 14648 34140 14724 34174
rect 14643 34117 14724 34140
rect 14539 34102 14724 34117
rect 14539 34083 14614 34102
rect 14539 34049 14609 34083
rect 14648 34068 14724 34102
rect 14643 34049 14724 34068
rect 14539 34030 14724 34049
rect 14539 34015 14614 34030
rect 14539 33981 14609 34015
rect 14648 33996 14724 34030
rect 14643 33981 14724 33996
rect 14539 33958 14724 33981
rect 14539 33947 14614 33958
rect 14539 33913 14609 33947
rect 14648 33924 14724 33958
rect 14643 33913 14724 33924
rect 14539 33886 14724 33913
rect 14539 33879 14614 33886
rect 14539 33845 14609 33879
rect 14648 33852 14724 33886
rect 14643 33845 14724 33852
rect 14539 33814 14724 33845
rect 14539 33811 14614 33814
rect 14539 33777 14609 33811
rect 14648 33780 14724 33814
rect 14643 33777 14724 33780
rect 14539 33743 14724 33777
rect 14539 33709 14609 33743
rect 14643 33742 14724 33743
rect 14539 33708 14614 33709
rect 14648 33708 14724 33742
rect 14539 33675 14724 33708
rect 14539 33641 14609 33675
rect 14643 33670 14724 33675
rect 14539 33636 14614 33641
rect 14648 33636 14724 33670
rect 14539 33607 14724 33636
rect 14539 33573 14609 33607
rect 14643 33598 14724 33607
rect 14539 33564 14614 33573
rect 14648 33564 14724 33598
rect 14539 33539 14724 33564
rect 14539 33505 14609 33539
rect 14643 33526 14724 33539
rect 14539 33492 14614 33505
rect 14648 33492 14724 33526
rect 14539 33471 14724 33492
rect 14539 33437 14609 33471
rect 14643 33454 14724 33471
rect 14539 33420 14614 33437
rect 14648 33420 14724 33454
rect 14539 33403 14724 33420
rect 14539 33369 14609 33403
rect 14643 33382 14724 33403
rect 14539 33348 14614 33369
rect 14648 33348 14724 33382
rect 14539 33335 14724 33348
rect 14539 33301 14609 33335
rect 14643 33310 14724 33335
rect 14539 33276 14614 33301
rect 14648 33276 14724 33310
rect 14539 33267 14724 33276
rect 14539 33233 14609 33267
rect 14643 33238 14724 33267
rect 14539 33204 14614 33233
rect 14648 33204 14724 33238
rect 14539 33199 14724 33204
rect 14539 33165 14609 33199
rect 14643 33166 14724 33199
rect 14539 33132 14614 33165
rect 14648 33132 14724 33166
rect 14539 33131 14724 33132
rect 14539 33097 14609 33131
rect 14643 33097 14724 33131
rect 14539 33094 14724 33097
rect 14539 33063 14614 33094
rect 14539 33029 14609 33063
rect 14648 33060 14724 33094
rect 14643 33029 14724 33060
rect 14539 33022 14724 33029
rect 14539 32995 14614 33022
rect 14539 32961 14609 32995
rect 14648 32988 14724 33022
rect 14643 32961 14724 32988
rect 14539 32950 14724 32961
rect 14539 32927 14614 32950
rect 14539 32893 14609 32927
rect 14648 32916 14724 32950
rect 14643 32893 14724 32916
rect 14539 32878 14724 32893
rect 14539 32859 14614 32878
rect 14539 32825 14609 32859
rect 14648 32844 14724 32878
rect 14643 32825 14724 32844
rect 14539 32806 14724 32825
rect 14539 32791 14614 32806
rect 14539 32757 14609 32791
rect 14648 32772 14724 32806
rect 14643 32757 14724 32772
rect 14539 32734 14724 32757
rect 14539 32723 14614 32734
rect 14539 32689 14609 32723
rect 14648 32700 14724 32734
rect 14643 32689 14724 32700
rect 14539 32662 14724 32689
rect 14539 32655 14614 32662
rect 14539 32621 14609 32655
rect 14648 32628 14724 32662
rect 14643 32621 14724 32628
rect 14539 32590 14724 32621
rect 14539 32587 14614 32590
rect 14539 32553 14609 32587
rect 14648 32556 14724 32590
rect 14643 32553 14724 32556
rect 14539 32519 14724 32553
rect 14539 32485 14609 32519
rect 14643 32518 14724 32519
rect 14539 32484 14614 32485
rect 14648 32484 14724 32518
rect 14539 32451 14724 32484
rect 14539 32417 14609 32451
rect 14643 32446 14724 32451
rect 14539 32412 14614 32417
rect 14648 32412 14724 32446
rect 14539 32383 14724 32412
rect 14539 32349 14609 32383
rect 14643 32374 14724 32383
rect 14539 32340 14614 32349
rect 14648 32340 14724 32374
rect 14539 32315 14724 32340
rect 14539 32281 14609 32315
rect 14643 32302 14724 32315
rect 14539 32268 14614 32281
rect 14648 32268 14724 32302
rect 14539 32247 14724 32268
rect 14539 32213 14609 32247
rect 14643 32230 14724 32247
rect 14539 32196 14614 32213
rect 14648 32196 14724 32230
rect 14539 32179 14724 32196
rect 14539 32145 14609 32179
rect 14643 32158 14724 32179
rect 14539 32124 14614 32145
rect 14648 32124 14724 32158
rect 14539 32111 14724 32124
rect 14539 32077 14609 32111
rect 14643 32086 14724 32111
rect 14539 32052 14614 32077
rect 14648 32052 14724 32086
rect 14539 32043 14724 32052
rect 14539 32009 14609 32043
rect 14643 32014 14724 32043
rect 14539 31980 14614 32009
rect 14648 31980 14724 32014
rect 14539 31975 14724 31980
rect 14539 31941 14609 31975
rect 14643 31942 14724 31975
rect 14539 31908 14614 31941
rect 14648 31908 14724 31942
rect 14539 31907 14724 31908
rect 14539 31873 14609 31907
rect 14643 31873 14724 31907
rect 14539 31870 14724 31873
rect 14539 31839 14614 31870
rect 14539 31805 14609 31839
rect 14648 31836 14724 31870
rect 14643 31805 14724 31836
rect 14539 31798 14724 31805
rect 14539 31771 14614 31798
rect 14539 31737 14609 31771
rect 14648 31764 14724 31798
rect 14643 31737 14724 31764
rect 14539 31726 14724 31737
rect 14539 31703 14614 31726
rect 14539 31669 14609 31703
rect 14648 31692 14724 31726
rect 14643 31669 14724 31692
rect 14539 31654 14724 31669
rect 14539 31635 14614 31654
rect 14539 31601 14609 31635
rect 14648 31620 14724 31654
rect 14643 31601 14724 31620
rect 14539 31582 14724 31601
rect 14539 31567 14614 31582
rect 14539 31533 14609 31567
rect 14648 31548 14724 31582
rect 14643 31533 14724 31548
rect 14539 31510 14724 31533
rect 14539 31499 14614 31510
rect 14539 31465 14609 31499
rect 14648 31476 14724 31510
rect 14643 31465 14724 31476
rect 14539 31438 14724 31465
rect 14539 31431 14614 31438
rect 14539 31397 14609 31431
rect 14648 31404 14724 31438
rect 14643 31397 14724 31404
rect 14539 31366 14724 31397
rect 14539 31363 14614 31366
rect 14539 31329 14609 31363
rect 14648 31332 14724 31366
rect 14643 31329 14724 31332
rect 14539 31295 14724 31329
rect 14539 31261 14609 31295
rect 14643 31294 14724 31295
rect 14539 31260 14614 31261
rect 14648 31260 14724 31294
rect 14539 31227 14724 31260
rect 14539 31193 14609 31227
rect 14643 31222 14724 31227
rect 14539 31188 14614 31193
rect 14648 31188 14724 31222
rect 14539 31159 14724 31188
rect 14539 31125 14609 31159
rect 14643 31150 14724 31159
rect 14539 31116 14614 31125
rect 14648 31116 14724 31150
rect 14539 31091 14724 31116
rect 14539 31057 14609 31091
rect 14643 31078 14724 31091
rect 14539 31044 14614 31057
rect 14648 31044 14724 31078
rect 14539 31023 14724 31044
rect 14539 30989 14609 31023
rect 14643 31006 14724 31023
rect 14539 30972 14614 30989
rect 14648 30972 14724 31006
rect 14539 30955 14724 30972
rect 14539 30921 14609 30955
rect 14643 30934 14724 30955
rect 14539 30900 14614 30921
rect 14648 30900 14724 30934
rect 14539 30887 14724 30900
rect 14539 30853 14609 30887
rect 14643 30862 14724 30887
rect 14539 30828 14614 30853
rect 14648 30828 14724 30862
rect 14539 30819 14724 30828
rect 14539 30785 14609 30819
rect 14643 30790 14724 30819
rect 14539 30756 14614 30785
rect 14648 30756 14724 30790
rect 14539 30751 14724 30756
rect 14539 30717 14609 30751
rect 14643 30718 14724 30751
rect 14539 30684 14614 30717
rect 14648 30684 14724 30718
rect 14539 30683 14724 30684
rect 14539 30649 14609 30683
rect 14643 30649 14724 30683
rect 14539 30646 14724 30649
rect 14539 30615 14614 30646
rect 14539 30581 14609 30615
rect 14648 30612 14724 30646
rect 14643 30581 14724 30612
rect 14539 30574 14724 30581
rect 14539 30547 14614 30574
rect 14539 30513 14609 30547
rect 14648 30540 14724 30574
rect 14643 30513 14724 30540
rect 14539 30502 14724 30513
rect 14539 30479 14614 30502
rect 14539 30445 14609 30479
rect 14648 30468 14724 30502
rect 14643 30445 14724 30468
rect 14539 30430 14724 30445
rect 14539 30411 14614 30430
rect 14539 30377 14609 30411
rect 14648 30396 14724 30430
rect 14643 30377 14724 30396
rect 14539 30358 14724 30377
rect 14539 30343 14614 30358
rect 14539 30309 14609 30343
rect 14648 30324 14724 30358
rect 14643 30309 14724 30324
rect 14539 30286 14724 30309
rect 14539 30275 14614 30286
rect 14539 30241 14609 30275
rect 14648 30252 14724 30286
rect 14643 30241 14724 30252
rect 14539 30214 14724 30241
rect 14539 30207 14614 30214
rect 14539 30173 14609 30207
rect 14648 30180 14724 30214
rect 14643 30173 14724 30180
rect 14539 30142 14724 30173
rect 14539 30139 14614 30142
rect 14539 30105 14609 30139
rect 14648 30108 14724 30142
rect 14643 30105 14724 30108
rect 14539 30071 14724 30105
rect 14539 30037 14609 30071
rect 14643 30070 14724 30071
rect 14539 30036 14614 30037
rect 14648 30036 14724 30070
rect 14539 30003 14724 30036
rect 14539 29969 14609 30003
rect 14643 29998 14724 30003
rect 14539 29964 14614 29969
rect 14648 29964 14724 29998
rect 14539 29935 14724 29964
rect 14539 29901 14609 29935
rect 14643 29926 14724 29935
rect 14539 29892 14614 29901
rect 14648 29892 14724 29926
rect 14539 29867 14724 29892
rect 14539 29833 14609 29867
rect 14643 29854 14724 29867
rect 14539 29820 14614 29833
rect 14648 29820 14724 29854
rect 14539 29799 14724 29820
rect 14539 29765 14609 29799
rect 14643 29782 14724 29799
rect 14539 29748 14614 29765
rect 14648 29748 14724 29782
rect 14539 29731 14724 29748
rect 14539 29697 14609 29731
rect 14643 29710 14724 29731
rect 14539 29676 14614 29697
rect 14648 29676 14724 29710
rect 14539 29663 14724 29676
rect 14539 29629 14609 29663
rect 14643 29638 14724 29663
rect 14539 29604 14614 29629
rect 14648 29604 14724 29638
rect 14539 29595 14724 29604
rect 14539 29561 14609 29595
rect 14643 29566 14724 29595
rect 14539 29532 14614 29561
rect 14648 29532 14724 29566
rect 14539 29527 14724 29532
rect 14539 29493 14609 29527
rect 14643 29494 14724 29527
rect 14539 29460 14614 29493
rect 14648 29460 14724 29494
rect 14539 29459 14724 29460
rect 14539 29425 14609 29459
rect 14643 29425 14724 29459
rect 14539 29422 14724 29425
rect 14539 29391 14614 29422
rect 14539 29357 14609 29391
rect 14648 29388 14724 29422
rect 14643 29357 14724 29388
rect 14539 29350 14724 29357
rect 14539 29323 14614 29350
rect 14539 29289 14609 29323
rect 14648 29316 14724 29350
rect 14643 29289 14724 29316
rect 14539 29278 14724 29289
rect 14539 29255 14614 29278
rect 14539 29221 14609 29255
rect 14648 29244 14724 29278
rect 14643 29221 14724 29244
rect 14539 29206 14724 29221
rect 14539 29187 14614 29206
rect 14539 29153 14609 29187
rect 14648 29172 14724 29206
rect 14643 29153 14724 29172
rect 14539 29134 14724 29153
rect 14539 29119 14614 29134
rect 14539 29085 14609 29119
rect 14648 29100 14724 29134
rect 14643 29085 14724 29100
rect 14539 29062 14724 29085
rect 14539 29051 14614 29062
rect 14539 29017 14609 29051
rect 14648 29028 14724 29062
rect 14643 29017 14724 29028
rect 14539 28990 14724 29017
rect 14539 28983 14614 28990
rect 14539 28949 14609 28983
rect 14648 28956 14724 28990
rect 14643 28949 14724 28956
rect 14539 28918 14724 28949
rect 14539 28915 14614 28918
rect 14539 28881 14609 28915
rect 14648 28884 14724 28918
rect 14643 28881 14724 28884
rect 14539 28847 14724 28881
rect 14539 28813 14609 28847
rect 14643 28846 14724 28847
rect 14539 28812 14614 28813
rect 14648 28812 14724 28846
rect 14539 28779 14724 28812
rect 14539 28745 14609 28779
rect 14643 28774 14724 28779
rect 14539 28740 14614 28745
rect 14648 28740 14724 28774
rect 14539 28711 14724 28740
rect 14539 28677 14609 28711
rect 14643 28702 14724 28711
rect 14539 28668 14614 28677
rect 14648 28668 14724 28702
rect 14539 28643 14724 28668
rect 14539 28609 14609 28643
rect 14643 28630 14724 28643
rect 14539 28596 14614 28609
rect 14648 28596 14724 28630
rect 14539 28575 14724 28596
rect 14539 28541 14609 28575
rect 14643 28558 14724 28575
rect 14539 28524 14614 28541
rect 14648 28524 14724 28558
rect 14539 28507 14724 28524
rect 14539 28473 14609 28507
rect 14643 28486 14724 28507
rect 14539 28452 14614 28473
rect 14648 28452 14724 28486
rect 14539 28439 14724 28452
rect 14539 28405 14609 28439
rect 14643 28414 14724 28439
rect 14539 28380 14614 28405
rect 14648 28380 14724 28414
rect 14539 28371 14724 28380
rect 14539 28337 14609 28371
rect 14643 28342 14724 28371
rect 14539 28308 14614 28337
rect 14648 28308 14724 28342
rect 14539 28303 14724 28308
rect 14539 28269 14609 28303
rect 14643 28270 14724 28303
rect 14539 28236 14614 28269
rect 14648 28236 14724 28270
rect 14539 28235 14724 28236
rect 14539 28201 14609 28235
rect 14643 28201 14724 28235
rect 14539 28198 14724 28201
rect 14539 28167 14614 28198
rect 14539 28133 14609 28167
rect 14648 28164 14724 28198
rect 14643 28133 14724 28164
rect 14539 28126 14724 28133
rect 14539 28099 14614 28126
rect 14539 28065 14609 28099
rect 14648 28092 14724 28126
rect 14643 28065 14724 28092
rect 14539 28054 14724 28065
rect 14539 28031 14614 28054
rect 14539 27997 14609 28031
rect 14648 28020 14724 28054
rect 14643 27997 14724 28020
rect 14539 27982 14724 27997
rect 14539 27963 14614 27982
rect 14539 27929 14609 27963
rect 14648 27948 14724 27982
rect 14643 27929 14724 27948
rect 14539 27910 14724 27929
rect 14539 27895 14614 27910
rect 14539 27861 14609 27895
rect 14648 27876 14724 27910
rect 14643 27861 14724 27876
rect 14539 27838 14724 27861
rect 14539 27827 14614 27838
rect 14539 27793 14609 27827
rect 14648 27804 14724 27838
rect 14643 27793 14724 27804
rect 14539 27766 14724 27793
rect 14539 27759 14614 27766
rect 14539 27725 14609 27759
rect 14648 27732 14724 27766
rect 14643 27725 14724 27732
rect 14539 27694 14724 27725
rect 14539 27691 14614 27694
rect 14539 27657 14609 27691
rect 14648 27660 14724 27694
rect 14643 27657 14724 27660
rect 14539 27623 14724 27657
rect 14539 27589 14609 27623
rect 14643 27622 14724 27623
rect 14539 27588 14614 27589
rect 14648 27588 14724 27622
rect 14539 27555 14724 27588
rect 14539 27521 14609 27555
rect 14643 27550 14724 27555
rect 14539 27516 14614 27521
rect 14648 27516 14724 27550
rect 14539 27487 14724 27516
rect 14539 27453 14609 27487
rect 14643 27478 14724 27487
rect 14539 27444 14614 27453
rect 14648 27444 14724 27478
rect 14539 27419 14724 27444
rect 14539 27385 14609 27419
rect 14643 27406 14724 27419
rect 14539 27372 14614 27385
rect 14648 27372 14724 27406
rect 14539 27351 14724 27372
rect 14539 27317 14609 27351
rect 14643 27334 14724 27351
rect 14539 27300 14614 27317
rect 14648 27300 14724 27334
rect 14539 27283 14724 27300
rect 14539 27249 14609 27283
rect 14643 27262 14724 27283
rect 14539 27228 14614 27249
rect 14648 27228 14724 27262
rect 14539 27215 14724 27228
rect 14539 27181 14609 27215
rect 14643 27190 14724 27215
rect 14539 27156 14614 27181
rect 14648 27156 14724 27190
rect 14539 27147 14724 27156
rect 14539 27113 14609 27147
rect 14643 27118 14724 27147
rect 14539 27084 14614 27113
rect 14648 27084 14724 27118
rect 14539 27079 14724 27084
rect 14539 27045 14609 27079
rect 14643 27046 14724 27079
rect 14539 27012 14614 27045
rect 14648 27012 14724 27046
rect 14539 27011 14724 27012
rect 14539 26977 14609 27011
rect 14643 26977 14724 27011
rect 14539 26974 14724 26977
rect 14539 26943 14614 26974
rect 14539 26909 14609 26943
rect 14648 26940 14724 26974
rect 14643 26909 14724 26940
rect 14539 26902 14724 26909
rect 14539 26875 14614 26902
rect 14539 26841 14609 26875
rect 14648 26868 14724 26902
rect 14643 26841 14724 26868
rect 14539 26830 14724 26841
rect 14539 26807 14614 26830
rect 14539 26773 14609 26807
rect 14648 26796 14724 26830
rect 14643 26773 14724 26796
rect 14539 26758 14724 26773
rect 14539 26739 14614 26758
rect 14539 26705 14609 26739
rect 14648 26724 14724 26758
rect 14643 26705 14724 26724
rect 14539 26686 14724 26705
rect 14539 26671 14614 26686
rect 14539 26637 14609 26671
rect 14648 26652 14724 26686
rect 14643 26637 14724 26652
rect 14539 26614 14724 26637
rect 14539 26603 14614 26614
rect 14539 26569 14609 26603
rect 14648 26580 14724 26614
rect 14643 26569 14724 26580
rect 14539 26542 14724 26569
rect 14539 26535 14614 26542
rect 14539 26501 14609 26535
rect 14648 26508 14724 26542
rect 14643 26501 14724 26508
rect 14539 26470 14724 26501
rect 14539 26467 14614 26470
rect 14539 26433 14609 26467
rect 14648 26436 14724 26470
rect 14643 26433 14724 26436
rect 14539 26399 14724 26433
rect 14539 26365 14609 26399
rect 14643 26398 14724 26399
rect 14539 26364 14614 26365
rect 14648 26364 14724 26398
rect 14539 26331 14724 26364
rect 14539 26297 14609 26331
rect 14643 26326 14724 26331
rect 14539 26292 14614 26297
rect 14648 26292 14724 26326
rect 14539 26263 14724 26292
rect 14539 26229 14609 26263
rect 14643 26254 14724 26263
rect 14539 26220 14614 26229
rect 14648 26220 14724 26254
rect 14539 26195 14724 26220
rect 14539 26161 14609 26195
rect 14643 26182 14724 26195
rect 14539 26148 14614 26161
rect 14648 26148 14724 26182
rect 14539 26127 14724 26148
rect 14539 26093 14609 26127
rect 14643 26110 14724 26127
rect 14539 26076 14614 26093
rect 14648 26076 14724 26110
rect 14539 26059 14724 26076
rect 14539 26025 14609 26059
rect 14643 26038 14724 26059
rect 14539 26004 14614 26025
rect 14648 26004 14724 26038
rect 14539 25991 14724 26004
rect 14539 25957 14609 25991
rect 14643 25966 14724 25991
rect 14539 25932 14614 25957
rect 14648 25932 14724 25966
rect 14539 25923 14724 25932
rect 14539 25889 14609 25923
rect 14643 25894 14724 25923
rect 14539 25860 14614 25889
rect 14648 25860 14724 25894
rect 14539 25855 14724 25860
rect 14539 25821 14609 25855
rect 14643 25822 14724 25855
rect 14539 25788 14614 25821
rect 14648 25788 14724 25822
rect 14539 25787 14724 25788
rect 14539 25753 14609 25787
rect 14643 25753 14724 25787
rect 14539 25750 14724 25753
rect 14539 25719 14614 25750
rect 14539 25685 14609 25719
rect 14648 25716 14724 25750
rect 14643 25685 14724 25716
rect 14539 25678 14724 25685
rect 14539 25651 14614 25678
rect 14539 25617 14609 25651
rect 14648 25644 14724 25678
rect 14643 25617 14724 25644
rect 14539 25606 14724 25617
rect 14539 25583 14614 25606
rect 14539 25549 14609 25583
rect 14648 25572 14724 25606
rect 14643 25549 14724 25572
rect 14539 25534 14724 25549
rect 14539 25515 14614 25534
rect 14539 25481 14609 25515
rect 14648 25500 14724 25534
rect 14643 25481 14724 25500
rect 14539 25462 14724 25481
rect 14539 25447 14614 25462
rect 14539 25413 14609 25447
rect 14648 25428 14724 25462
rect 14643 25413 14724 25428
rect 14539 25390 14724 25413
rect 14539 25379 14614 25390
rect 14539 25345 14609 25379
rect 14648 25356 14724 25390
rect 14643 25345 14724 25356
rect 14539 25318 14724 25345
rect 14539 25311 14614 25318
rect 14539 25277 14609 25311
rect 14648 25284 14724 25318
rect 14643 25277 14724 25284
rect 14539 25246 14724 25277
rect 14539 25243 14614 25246
rect 14539 25209 14609 25243
rect 14648 25212 14724 25246
rect 14643 25209 14724 25212
rect 14539 25175 14724 25209
rect 14539 25141 14609 25175
rect 14643 25174 14724 25175
rect 14539 25140 14614 25141
rect 14648 25140 14724 25174
rect 14539 25107 14724 25140
rect 14539 25073 14609 25107
rect 14643 25102 14724 25107
rect 14539 25068 14614 25073
rect 14648 25068 14724 25102
rect 14539 25039 14724 25068
rect 14539 25005 14609 25039
rect 14643 25030 14724 25039
rect 14539 24996 14614 25005
rect 14648 24996 14724 25030
rect 14539 24971 14724 24996
rect 14539 24937 14609 24971
rect 14643 24958 14724 24971
rect 14539 24924 14614 24937
rect 14648 24924 14724 24958
rect 14539 24903 14724 24924
rect 14539 24869 14609 24903
rect 14643 24886 14724 24903
rect 14539 24852 14614 24869
rect 14648 24852 14724 24886
rect 14539 24835 14724 24852
rect 14539 24801 14609 24835
rect 14643 24814 14724 24835
rect 14539 24780 14614 24801
rect 14648 24780 14724 24814
rect 14539 24767 14724 24780
rect 14539 24733 14609 24767
rect 14643 24742 14724 24767
rect 14539 24708 14614 24733
rect 14648 24708 14724 24742
rect 14539 24699 14724 24708
rect 14539 24665 14609 24699
rect 14643 24670 14724 24699
rect 14539 24636 14614 24665
rect 14648 24636 14724 24670
rect 14539 24631 14724 24636
rect 14539 24597 14609 24631
rect 14643 24598 14724 24631
rect 14539 24564 14614 24597
rect 14648 24564 14724 24598
rect 14539 24563 14724 24564
rect 14539 24529 14609 24563
rect 14643 24529 14724 24563
rect 14539 24526 14724 24529
rect 14539 24495 14614 24526
rect 14539 24461 14609 24495
rect 14648 24492 14724 24526
rect 14643 24461 14724 24492
rect 14539 24454 14724 24461
rect 14539 24427 14614 24454
rect 14539 24393 14609 24427
rect 14648 24420 14724 24454
rect 14643 24393 14724 24420
rect 14539 24382 14724 24393
rect 14539 24359 14614 24382
rect 14539 24325 14609 24359
rect 14648 24348 14724 24382
rect 14643 24325 14724 24348
rect 14539 24310 14724 24325
rect 14539 24291 14614 24310
rect 14539 24257 14609 24291
rect 14648 24276 14724 24310
rect 14643 24257 14724 24276
rect 14539 24238 14724 24257
rect 14539 24223 14614 24238
rect 14539 24189 14609 24223
rect 14648 24204 14724 24238
rect 14643 24189 14724 24204
rect 14539 24166 14724 24189
rect 14539 24155 14614 24166
rect 14539 24121 14609 24155
rect 14648 24132 14724 24166
rect 14643 24121 14724 24132
rect 14539 24094 14724 24121
rect 14539 24087 14614 24094
rect 14539 24053 14609 24087
rect 14648 24060 14724 24094
rect 14643 24053 14724 24060
rect 14539 24022 14724 24053
rect 14539 24019 14614 24022
rect 14539 23985 14609 24019
rect 14648 23988 14724 24022
rect 14643 23985 14724 23988
rect 14539 23951 14724 23985
rect 14539 23917 14609 23951
rect 14643 23950 14724 23951
rect 14539 23916 14614 23917
rect 14648 23916 14724 23950
rect 14539 23883 14724 23916
rect 14539 23849 14609 23883
rect 14643 23878 14724 23883
rect 14539 23844 14614 23849
rect 14648 23844 14724 23878
rect 14539 23815 14724 23844
rect 14539 23781 14609 23815
rect 14643 23806 14724 23815
rect 14539 23772 14614 23781
rect 14648 23772 14724 23806
rect 14539 23747 14724 23772
rect 14539 23713 14609 23747
rect 14643 23734 14724 23747
rect 14539 23700 14614 23713
rect 14648 23700 14724 23734
rect 14539 23679 14724 23700
rect 14539 23645 14609 23679
rect 14643 23662 14724 23679
rect 14539 23628 14614 23645
rect 14648 23628 14724 23662
rect 14539 23611 14724 23628
rect 14539 23577 14609 23611
rect 14643 23590 14724 23611
rect 14539 23556 14614 23577
rect 14648 23556 14724 23590
rect 14539 23543 14724 23556
rect 14539 23509 14609 23543
rect 14643 23518 14724 23543
rect 14539 23484 14614 23509
rect 14648 23484 14724 23518
rect 14539 23475 14724 23484
rect 14539 23441 14609 23475
rect 14643 23446 14724 23475
rect 14539 23412 14614 23441
rect 14648 23412 14724 23446
rect 14539 23407 14724 23412
rect 14539 23373 14609 23407
rect 14643 23374 14724 23407
rect 14539 23340 14614 23373
rect 14648 23340 14724 23374
rect 14539 23339 14724 23340
rect 14539 23305 14609 23339
rect 14643 23305 14724 23339
rect 14539 23302 14724 23305
rect 14539 23271 14614 23302
rect 14539 23237 14609 23271
rect 14648 23268 14724 23302
rect 14643 23237 14724 23268
rect 14539 23230 14724 23237
rect 14539 23203 14614 23230
rect 14539 23169 14609 23203
rect 14648 23196 14724 23230
rect 14643 23169 14724 23196
rect 14539 23158 14724 23169
rect 14539 23135 14614 23158
rect 14539 23101 14609 23135
rect 14648 23124 14724 23158
rect 14643 23101 14724 23124
rect 14539 23086 14724 23101
rect 14539 23067 14614 23086
rect 14539 23033 14609 23067
rect 14648 23052 14724 23086
rect 14643 23033 14724 23052
rect 14539 23014 14724 23033
rect 14539 22999 14614 23014
rect 14539 22965 14609 22999
rect 14648 22980 14724 23014
rect 14643 22965 14724 22980
rect 14539 22942 14724 22965
rect 14539 22931 14614 22942
rect 14539 22897 14609 22931
rect 14648 22908 14724 22942
rect 14643 22897 14724 22908
rect 14539 22870 14724 22897
rect 14539 22863 14614 22870
rect 14539 22829 14609 22863
rect 14648 22836 14724 22870
rect 14643 22829 14724 22836
rect 14539 22798 14724 22829
rect 14539 22795 14614 22798
rect 14539 22761 14609 22795
rect 14648 22764 14724 22798
rect 14643 22761 14724 22764
rect 14539 22727 14724 22761
rect 14539 22693 14609 22727
rect 14643 22726 14724 22727
rect 14539 22692 14614 22693
rect 14648 22692 14724 22726
rect 14539 22659 14724 22692
rect 14539 22625 14609 22659
rect 14643 22654 14724 22659
rect 14539 22620 14614 22625
rect 14648 22620 14724 22654
rect 14539 22591 14724 22620
rect 14539 22557 14609 22591
rect 14643 22582 14724 22591
rect 14539 22548 14614 22557
rect 14648 22548 14724 22582
rect 14539 22523 14724 22548
rect 14539 22489 14609 22523
rect 14643 22510 14724 22523
rect 14539 22476 14614 22489
rect 14648 22476 14724 22510
rect 14539 22455 14724 22476
rect 14539 22421 14609 22455
rect 14643 22438 14724 22455
rect 14539 22404 14614 22421
rect 14648 22404 14724 22438
rect 14539 22387 14724 22404
rect 14539 22353 14609 22387
rect 14643 22366 14724 22387
rect 14539 22332 14614 22353
rect 14648 22332 14724 22366
rect 14539 22319 14724 22332
rect 14539 22285 14609 22319
rect 14643 22294 14724 22319
rect 14539 22260 14614 22285
rect 14648 22260 14724 22294
rect 14539 22251 14724 22260
rect 14539 22217 14609 22251
rect 14643 22222 14724 22251
rect 14539 22188 14614 22217
rect 14648 22188 14724 22222
rect 14539 22183 14724 22188
rect 14539 22149 14609 22183
rect 14643 22150 14724 22183
rect 14539 22116 14614 22149
rect 14648 22116 14724 22150
rect 14539 22115 14724 22116
rect 14539 22081 14609 22115
rect 14643 22081 14724 22115
rect 14539 22078 14724 22081
rect 14539 22047 14614 22078
rect 14539 22013 14609 22047
rect 14648 22044 14724 22078
rect 14643 22013 14724 22044
rect 14539 22006 14724 22013
rect 14539 21979 14614 22006
rect 14539 21945 14609 21979
rect 14648 21972 14724 22006
rect 14643 21945 14724 21972
rect 14539 21934 14724 21945
rect 14539 21911 14614 21934
rect 14539 21877 14609 21911
rect 14648 21900 14724 21934
rect 14643 21877 14724 21900
rect 14539 21862 14724 21877
rect 14539 21843 14614 21862
rect 14539 21809 14609 21843
rect 14648 21828 14724 21862
rect 14643 21809 14724 21828
rect 14539 21790 14724 21809
rect 14539 21775 14614 21790
rect 14539 21741 14609 21775
rect 14648 21756 14724 21790
rect 14643 21741 14724 21756
rect 14539 21718 14724 21741
rect 14539 21707 14614 21718
rect 14539 21673 14609 21707
rect 14648 21684 14724 21718
rect 14643 21673 14724 21684
rect 14539 21646 14724 21673
rect 14539 21639 14614 21646
rect 14539 21605 14609 21639
rect 14648 21612 14724 21646
rect 14643 21605 14724 21612
rect 14539 21574 14724 21605
rect 14539 21571 14614 21574
rect 14539 21537 14609 21571
rect 14648 21540 14724 21574
rect 14643 21537 14724 21540
rect 14539 21503 14724 21537
rect 14539 21469 14609 21503
rect 14643 21502 14724 21503
rect 14539 21468 14614 21469
rect 14648 21468 14724 21502
rect 14539 21435 14724 21468
rect 14539 21401 14609 21435
rect 14643 21430 14724 21435
rect 14539 21396 14614 21401
rect 14648 21396 14724 21430
rect 14539 21367 14724 21396
rect 14539 21333 14609 21367
rect 14643 21358 14724 21367
rect 14539 21324 14614 21333
rect 14648 21324 14724 21358
rect 14539 21299 14724 21324
rect 14539 21265 14609 21299
rect 14643 21286 14724 21299
rect 14539 21252 14614 21265
rect 14648 21252 14724 21286
rect 14539 21231 14724 21252
rect 14539 21197 14609 21231
rect 14643 21214 14724 21231
rect 14539 21180 14614 21197
rect 14648 21180 14724 21214
rect 14539 21163 14724 21180
rect 14539 21129 14609 21163
rect 14643 21142 14724 21163
rect 14539 21108 14614 21129
rect 14648 21108 14724 21142
rect 14539 21095 14724 21108
rect 14539 21061 14609 21095
rect 14643 21070 14724 21095
rect 14539 21036 14614 21061
rect 14648 21036 14724 21070
rect 14539 21027 14724 21036
rect 14539 20993 14609 21027
rect 14643 20998 14724 21027
rect 14539 20964 14614 20993
rect 14648 20964 14724 20998
rect 14539 20959 14724 20964
rect 14539 20925 14609 20959
rect 14643 20926 14724 20959
rect 14539 20892 14614 20925
rect 14648 20892 14724 20926
rect 14539 20891 14724 20892
rect 14539 20857 14609 20891
rect 14643 20857 14724 20891
rect 14539 20854 14724 20857
rect 14539 20823 14614 20854
rect 14539 20789 14609 20823
rect 14648 20820 14724 20854
rect 14643 20789 14724 20820
rect 14539 20782 14724 20789
rect 14539 20755 14614 20782
rect 14539 20721 14609 20755
rect 14648 20748 14724 20782
rect 14643 20721 14724 20748
rect 14539 20710 14724 20721
rect 14539 20687 14614 20710
rect 14539 20653 14609 20687
rect 14648 20676 14724 20710
rect 14643 20653 14724 20676
rect 14539 20638 14724 20653
rect 14539 20619 14614 20638
rect 14539 20585 14609 20619
rect 14648 20604 14724 20638
rect 14643 20585 14724 20604
rect 14539 20566 14724 20585
rect 14539 20551 14614 20566
rect 14539 20517 14609 20551
rect 14648 20532 14724 20566
rect 14643 20517 14724 20532
rect 14539 20494 14724 20517
rect 14539 20483 14614 20494
rect 14539 20449 14609 20483
rect 14648 20460 14724 20494
rect 14643 20449 14724 20460
rect 14539 20422 14724 20449
rect 14539 20415 14614 20422
rect 14539 20381 14609 20415
rect 14648 20388 14724 20422
rect 14643 20381 14724 20388
rect 14539 20350 14724 20381
rect 14539 20347 14614 20350
rect 14539 20313 14609 20347
rect 14648 20316 14724 20350
rect 14643 20313 14724 20316
rect 14539 20279 14724 20313
rect 14539 20245 14609 20279
rect 14643 20278 14724 20279
rect 14539 20244 14614 20245
rect 14648 20244 14724 20278
rect 14539 20211 14724 20244
rect 14539 20177 14609 20211
rect 14643 20206 14724 20211
rect 14539 20172 14614 20177
rect 14648 20172 14724 20206
rect 14539 20143 14724 20172
rect 14539 20109 14609 20143
rect 14643 20134 14724 20143
rect 14539 20100 14614 20109
rect 14648 20100 14724 20134
rect 14539 20075 14724 20100
rect 14539 20041 14609 20075
rect 14643 20062 14724 20075
rect 14539 20028 14614 20041
rect 14648 20028 14724 20062
rect 14539 20007 14724 20028
rect 14539 19973 14609 20007
rect 14643 19990 14724 20007
rect 14539 19956 14614 19973
rect 14648 19956 14724 19990
rect 14539 19939 14724 19956
rect 14539 19905 14609 19939
rect 14643 19918 14724 19939
rect 14539 19884 14614 19905
rect 14648 19884 14724 19918
rect 14539 19871 14724 19884
rect 14539 19837 14609 19871
rect 14643 19846 14724 19871
rect 14539 19812 14614 19837
rect 14648 19812 14724 19846
rect 14539 19803 14724 19812
rect 14539 19769 14609 19803
rect 14643 19774 14724 19803
rect 14539 19740 14614 19769
rect 14648 19740 14724 19774
rect 14539 19735 14724 19740
rect 14539 19701 14609 19735
rect 14643 19702 14724 19735
rect 14539 19668 14614 19701
rect 14648 19668 14724 19702
rect 14539 19667 14724 19668
rect 14539 19633 14609 19667
rect 14643 19633 14724 19667
rect 14539 19630 14724 19633
rect 14539 19599 14614 19630
rect 14539 19565 14609 19599
rect 14648 19596 14724 19630
rect 14643 19565 14724 19596
rect 14539 19558 14724 19565
rect 14539 19531 14614 19558
rect 14539 19497 14609 19531
rect 14648 19524 14724 19558
rect 14643 19497 14724 19524
rect 14539 19486 14724 19497
rect 14539 19463 14614 19486
rect 14539 19429 14609 19463
rect 14648 19452 14724 19486
rect 14643 19429 14724 19452
rect 14539 19414 14724 19429
rect 14539 19395 14614 19414
rect 14539 19361 14609 19395
rect 14648 19380 14724 19414
rect 14643 19361 14724 19380
rect 14539 19342 14724 19361
rect 14539 19327 14614 19342
rect 14539 19293 14609 19327
rect 14648 19308 14724 19342
rect 14643 19293 14724 19308
rect 14539 19270 14724 19293
rect 14539 19259 14614 19270
rect 14539 19225 14609 19259
rect 14648 19236 14724 19270
rect 14643 19225 14724 19236
rect 14539 19198 14724 19225
rect 14539 19191 14614 19198
rect 14539 19157 14609 19191
rect 14648 19164 14724 19198
rect 14643 19157 14724 19164
rect 14539 19126 14724 19157
rect 14539 19123 14614 19126
rect 14539 19089 14609 19123
rect 14648 19092 14724 19126
rect 14643 19089 14724 19092
rect 14539 19055 14724 19089
rect 14539 19021 14609 19055
rect 14643 19054 14724 19055
rect 14539 19020 14614 19021
rect 14648 19020 14724 19054
rect 14539 18987 14724 19020
rect 14539 18953 14609 18987
rect 14643 18982 14724 18987
rect 14539 18948 14614 18953
rect 14648 18948 14724 18982
rect 14539 18919 14724 18948
rect 14539 18885 14609 18919
rect 14643 18910 14724 18919
rect 14539 18876 14614 18885
rect 14648 18876 14724 18910
rect 14539 18851 14724 18876
rect 14539 18817 14609 18851
rect 14643 18838 14724 18851
rect 14539 18804 14614 18817
rect 14648 18804 14724 18838
rect 14539 18783 14724 18804
rect 14539 18749 14609 18783
rect 14643 18766 14724 18783
rect 14539 18732 14614 18749
rect 14648 18732 14724 18766
rect 14539 18715 14724 18732
rect 14539 18681 14609 18715
rect 14643 18694 14724 18715
rect 14539 18660 14614 18681
rect 14648 18660 14724 18694
rect 14539 18647 14724 18660
rect 14539 18613 14609 18647
rect 14643 18622 14724 18647
rect 14539 18588 14614 18613
rect 14648 18588 14724 18622
rect 14539 18579 14724 18588
rect 14539 18545 14609 18579
rect 14643 18550 14724 18579
rect 14539 18516 14614 18545
rect 14648 18516 14724 18550
rect 14539 18511 14724 18516
rect 14539 18477 14609 18511
rect 14643 18478 14724 18511
rect 14539 18444 14614 18477
rect 14648 18444 14724 18478
rect 14539 18443 14724 18444
rect 14539 18409 14609 18443
rect 14643 18409 14724 18443
rect 14539 18406 14724 18409
rect 14539 18375 14614 18406
rect 14539 18341 14609 18375
rect 14648 18372 14724 18406
rect 14643 18341 14724 18372
rect 14539 18334 14724 18341
rect 14539 18307 14614 18334
rect 14539 18273 14609 18307
rect 14648 18300 14724 18334
rect 14643 18273 14724 18300
rect 14539 18262 14724 18273
rect 14539 18239 14614 18262
rect 14539 18205 14609 18239
rect 14648 18228 14724 18262
rect 14643 18205 14724 18228
rect 14539 18190 14724 18205
rect 14539 18171 14614 18190
rect 14539 18137 14609 18171
rect 14648 18156 14724 18190
rect 14643 18137 14724 18156
rect 14539 18118 14724 18137
rect 14539 18103 14614 18118
rect 14539 18069 14609 18103
rect 14648 18084 14724 18118
rect 14643 18069 14724 18084
rect 14539 18046 14724 18069
rect 14539 18035 14614 18046
rect 14539 18001 14609 18035
rect 14648 18012 14724 18046
rect 14643 18001 14724 18012
rect 14539 17974 14724 18001
rect 14539 17967 14614 17974
rect 14539 17933 14609 17967
rect 14648 17940 14724 17974
rect 14643 17933 14724 17940
rect 14539 17902 14724 17933
rect 14539 17899 14614 17902
rect 14539 17865 14609 17899
rect 14648 17868 14724 17902
rect 14643 17865 14724 17868
rect 14539 17831 14724 17865
rect 14539 17797 14609 17831
rect 14643 17830 14724 17831
rect 14539 17796 14614 17797
rect 14648 17796 14724 17830
rect 14539 17763 14724 17796
rect 14539 17729 14609 17763
rect 14643 17758 14724 17763
rect 14539 17724 14614 17729
rect 14648 17724 14724 17758
rect 14539 17695 14724 17724
rect 14539 17661 14609 17695
rect 14643 17686 14724 17695
rect 14539 17652 14614 17661
rect 14648 17652 14724 17686
rect 14539 17627 14724 17652
rect 14539 17593 14609 17627
rect 14643 17614 14724 17627
rect 14539 17580 14614 17593
rect 14648 17580 14724 17614
rect 14539 17559 14724 17580
rect 14539 17525 14609 17559
rect 14643 17542 14724 17559
rect 14539 17508 14614 17525
rect 14648 17508 14724 17542
rect 14539 17491 14724 17508
rect 14539 17457 14609 17491
rect 14643 17470 14724 17491
rect 14539 17436 14614 17457
rect 14648 17436 14724 17470
rect 14539 17423 14724 17436
rect 14539 17389 14609 17423
rect 14643 17398 14724 17423
rect 14539 17364 14614 17389
rect 14648 17364 14724 17398
rect 14539 17355 14724 17364
rect 14539 17321 14609 17355
rect 14643 17326 14724 17355
rect 14539 17292 14614 17321
rect 14648 17292 14724 17326
rect 14539 17287 14724 17292
rect 14539 17253 14609 17287
rect 14643 17254 14724 17287
rect 14539 17220 14614 17253
rect 14648 17220 14724 17254
rect 14539 17219 14724 17220
rect 14539 17185 14609 17219
rect 14643 17185 14724 17219
rect 14539 17182 14724 17185
rect 14539 17151 14614 17182
rect 14539 17117 14609 17151
rect 14648 17148 14724 17182
rect 14643 17117 14724 17148
rect 14539 17110 14724 17117
rect 14539 17083 14614 17110
rect 14539 17049 14609 17083
rect 14648 17076 14724 17110
rect 14643 17049 14724 17076
rect 14539 17038 14724 17049
rect 14539 17015 14614 17038
rect 14539 16981 14609 17015
rect 14648 17004 14724 17038
rect 14643 16981 14724 17004
rect 14539 16966 14724 16981
rect 14539 16947 14614 16966
rect 14539 16913 14609 16947
rect 14648 16932 14724 16966
rect 14643 16913 14724 16932
rect 14539 16894 14724 16913
rect 14539 16879 14614 16894
rect 14539 16845 14609 16879
rect 14648 16860 14724 16894
rect 14643 16845 14724 16860
rect 14539 16822 14724 16845
rect 14539 16811 14614 16822
rect 14539 16777 14609 16811
rect 14648 16788 14724 16822
rect 14643 16777 14724 16788
rect 14539 16750 14724 16777
rect 14539 16743 14614 16750
rect 14539 16709 14609 16743
rect 14648 16716 14724 16750
rect 14643 16709 14724 16716
rect 14539 16678 14724 16709
rect 14539 16675 14614 16678
rect 14539 16641 14609 16675
rect 14648 16644 14724 16678
rect 14643 16641 14724 16644
rect 14539 16607 14724 16641
rect 14539 16573 14609 16607
rect 14643 16606 14724 16607
rect 14539 16572 14614 16573
rect 14648 16572 14724 16606
rect 14539 16539 14724 16572
rect 14539 16505 14609 16539
rect 14643 16534 14724 16539
rect 14539 16500 14614 16505
rect 14648 16500 14724 16534
rect 14539 16471 14724 16500
rect 14539 16437 14609 16471
rect 14643 16462 14724 16471
rect 14539 16428 14614 16437
rect 14648 16428 14724 16462
rect 14539 16403 14724 16428
rect 14539 16369 14609 16403
rect 14643 16390 14724 16403
rect 14539 16356 14614 16369
rect 14648 16356 14724 16390
rect 14539 16335 14724 16356
rect 14539 16301 14609 16335
rect 14643 16318 14724 16335
rect 14539 16284 14614 16301
rect 14648 16284 14724 16318
rect 14539 16267 14724 16284
rect 14539 16233 14609 16267
rect 14643 16246 14724 16267
rect 14539 16212 14614 16233
rect 14648 16212 14724 16246
rect 14539 16199 14724 16212
rect 14539 16165 14609 16199
rect 14643 16174 14724 16199
rect 14539 16140 14614 16165
rect 14648 16140 14724 16174
rect 14539 16131 14724 16140
rect 14539 16097 14609 16131
rect 14643 16102 14724 16131
rect 14539 16068 14614 16097
rect 14648 16068 14724 16102
rect 14539 16063 14724 16068
rect 14539 16029 14609 16063
rect 14643 16030 14724 16063
rect 14539 15996 14614 16029
rect 14648 15996 14724 16030
rect 14539 15995 14724 15996
rect 14539 15961 14609 15995
rect 14643 15961 14724 15995
rect 14539 15958 14724 15961
rect 14539 15927 14614 15958
rect 14539 15893 14609 15927
rect 14648 15924 14724 15958
rect 14643 15893 14724 15924
rect 14539 15886 14724 15893
rect 14539 15859 14614 15886
rect 14539 15825 14609 15859
rect 14648 15852 14724 15886
rect 14643 15825 14724 15852
rect 14539 15814 14724 15825
rect 14539 15791 14614 15814
rect 14539 15757 14609 15791
rect 14648 15780 14724 15814
rect 14643 15757 14724 15780
rect 14539 15742 14724 15757
rect 14539 15723 14614 15742
rect 14539 15689 14609 15723
rect 14648 15708 14724 15742
rect 14643 15689 14724 15708
rect 14539 15670 14724 15689
rect 14539 15655 14614 15670
rect 14539 15621 14609 15655
rect 14648 15636 14724 15670
rect 14643 15621 14724 15636
rect 14539 15598 14724 15621
rect 14539 15587 14614 15598
rect 14539 15553 14609 15587
rect 14648 15564 14724 15598
rect 14643 15553 14724 15564
rect 14539 15526 14724 15553
rect 14539 15519 14614 15526
rect 14539 15485 14609 15519
rect 14648 15492 14724 15526
rect 14643 15485 14724 15492
rect 14539 15454 14724 15485
rect 14539 15451 14614 15454
rect 14539 15417 14609 15451
rect 14648 15420 14724 15454
rect 14643 15417 14724 15420
rect 14539 15383 14724 15417
rect 14539 15349 14609 15383
rect 14643 15382 14724 15383
rect 14539 15348 14614 15349
rect 14648 15348 14724 15382
rect 14539 15315 14724 15348
rect 14539 15281 14609 15315
rect 14643 15310 14724 15315
rect 14539 15276 14614 15281
rect 14648 15276 14724 15310
rect 14539 15247 14724 15276
rect 14539 15213 14609 15247
rect 14643 15238 14724 15247
rect 14539 15204 14614 15213
rect 14648 15204 14724 15238
rect 14539 15179 14724 15204
rect 14539 15145 14609 15179
rect 14643 15166 14724 15179
rect 14539 15132 14614 15145
rect 14648 15132 14724 15166
rect 14539 15111 14724 15132
rect 14539 15077 14609 15111
rect 14643 15094 14724 15111
rect 14539 15060 14614 15077
rect 14648 15060 14724 15094
rect 14539 15043 14724 15060
rect 14539 15009 14609 15043
rect 14643 15022 14724 15043
rect 14539 14988 14614 15009
rect 14648 14988 14724 15022
rect 14539 14975 14724 14988
rect 14539 14941 14609 14975
rect 14643 14950 14724 14975
rect 14539 14916 14614 14941
rect 14648 14916 14724 14950
rect 14539 14907 14724 14916
rect 14539 14873 14609 14907
rect 14643 14878 14724 14907
rect 14539 14844 14614 14873
rect 14648 14844 14724 14878
rect 14539 14839 14724 14844
rect 14539 14805 14609 14839
rect 14643 14806 14724 14839
rect 14539 14772 14614 14805
rect 14648 14772 14724 14806
rect 14539 14771 14724 14772
rect 14539 14737 14609 14771
rect 14643 14737 14724 14771
rect 14539 14734 14724 14737
rect 14539 14703 14614 14734
rect 14539 14669 14609 14703
rect 14648 14700 14724 14734
rect 14643 14669 14724 14700
rect 14539 14662 14724 14669
rect 14539 14635 14614 14662
rect 14539 14601 14609 14635
rect 14648 14628 14724 14662
rect 14643 14601 14724 14628
rect 14539 14590 14724 14601
rect 14539 14567 14614 14590
rect 14539 14533 14609 14567
rect 14648 14556 14724 14590
rect 14643 14533 14724 14556
rect 14539 14518 14724 14533
rect 14539 14499 14614 14518
rect 14539 14465 14609 14499
rect 14648 14484 14724 14518
rect 14643 14465 14724 14484
rect 14539 14446 14724 14465
rect 14539 14431 14614 14446
rect 14539 14397 14609 14431
rect 14648 14412 14724 14446
rect 14643 14397 14724 14412
rect 14539 14374 14724 14397
rect 14539 14363 14614 14374
rect 14539 14329 14609 14363
rect 14648 14340 14724 14374
rect 14643 14329 14724 14340
rect 14539 14302 14724 14329
rect 14539 14295 14614 14302
rect 14539 14261 14609 14295
rect 14648 14268 14724 14302
rect 14643 14261 14724 14268
rect 14539 14230 14724 14261
rect 14539 14227 14614 14230
rect 14539 14193 14609 14227
rect 14648 14196 14724 14230
rect 14643 14193 14724 14196
rect 14539 14159 14724 14193
rect 14539 14125 14609 14159
rect 14643 14158 14724 14159
rect 14539 14124 14614 14125
rect 14648 14124 14724 14158
rect 14539 14091 14724 14124
rect 14539 14057 14609 14091
rect 14643 14086 14724 14091
rect 14539 14052 14614 14057
rect 14648 14052 14724 14086
rect 14539 14023 14724 14052
rect 14539 13989 14609 14023
rect 14643 14014 14724 14023
rect 14539 13980 14614 13989
rect 14648 13980 14724 14014
rect 14539 13955 14724 13980
rect 14539 13921 14609 13955
rect 14643 13942 14724 13955
rect 14539 13908 14614 13921
rect 14648 13908 14724 13942
rect 14539 13887 14724 13908
rect 14539 13853 14609 13887
rect 14643 13870 14724 13887
rect 14539 13836 14614 13853
rect 14648 13836 14724 13870
rect 14539 13819 14724 13836
rect 14539 13785 14609 13819
rect 14643 13798 14724 13819
rect 14539 13764 14614 13785
rect 14648 13764 14724 13798
rect 14539 13751 14724 13764
rect 14539 13717 14609 13751
rect 14643 13726 14724 13751
rect 14539 13692 14614 13717
rect 14648 13692 14724 13726
rect 14539 13683 14724 13692
rect 14539 13649 14609 13683
rect 14643 13654 14724 13683
rect 14539 13620 14614 13649
rect 14648 13620 14724 13654
rect 14539 13615 14724 13620
rect 14539 13581 14609 13615
rect 14643 13582 14724 13615
rect 14539 13548 14614 13581
rect 14648 13548 14724 13582
rect 14539 13547 14724 13548
rect 14539 13513 14609 13547
rect 14643 13513 14724 13547
rect 14539 13510 14724 13513
rect 14539 13479 14614 13510
rect 14539 13445 14609 13479
rect 14648 13476 14724 13510
rect 14643 13445 14724 13476
rect 14539 13438 14724 13445
rect 14539 13411 14614 13438
rect 14539 13377 14609 13411
rect 14648 13404 14724 13438
rect 14643 13377 14724 13404
rect 14539 13366 14724 13377
rect 14539 13343 14614 13366
rect 14539 13309 14609 13343
rect 14648 13332 14724 13366
rect 14643 13309 14724 13332
rect 14539 13294 14724 13309
rect 14539 13275 14614 13294
rect 14539 13241 14609 13275
rect 14648 13260 14724 13294
rect 14643 13241 14724 13260
rect 14539 13222 14724 13241
rect 14539 13207 14614 13222
rect 14539 13173 14609 13207
rect 14648 13188 14724 13222
rect 14643 13173 14724 13188
rect 14539 13150 14724 13173
rect 14539 13139 14614 13150
rect 14539 13105 14609 13139
rect 14648 13116 14724 13150
rect 14643 13105 14724 13116
rect 14539 13078 14724 13105
rect 14539 13071 14614 13078
rect 14539 13037 14609 13071
rect 14648 13044 14724 13078
rect 14643 13037 14724 13044
rect 14539 13006 14724 13037
rect 14539 13003 14614 13006
rect 14539 12969 14609 13003
rect 14648 12972 14724 13006
rect 14643 12969 14724 12972
rect 14539 12935 14724 12969
rect 14539 12901 14609 12935
rect 14643 12934 14724 12935
rect 14539 12900 14614 12901
rect 14648 12900 14724 12934
rect 14539 12867 14724 12900
rect 14539 12833 14609 12867
rect 14643 12862 14724 12867
rect 14539 12828 14614 12833
rect 14648 12828 14724 12862
rect 14539 12799 14724 12828
rect 14539 12765 14609 12799
rect 14643 12790 14724 12799
rect 14539 12756 14614 12765
rect 14648 12756 14724 12790
rect 14539 12731 14724 12756
rect 14539 12697 14609 12731
rect 14643 12718 14724 12731
rect 14539 12684 14614 12697
rect 14648 12684 14724 12718
rect 14539 12663 14724 12684
rect 14539 12629 14609 12663
rect 14643 12646 14724 12663
rect 14539 12612 14614 12629
rect 14648 12612 14724 12646
rect 14539 12595 14724 12612
rect 14539 12561 14609 12595
rect 14643 12574 14724 12595
rect 14539 12540 14614 12561
rect 14648 12540 14724 12574
rect 14539 12527 14724 12540
rect 14539 12493 14609 12527
rect 14643 12502 14724 12527
rect 14539 12468 14614 12493
rect 14648 12468 14724 12502
rect 14539 12459 14724 12468
rect 14539 12425 14609 12459
rect 14643 12430 14724 12459
rect 14539 12396 14614 12425
rect 14648 12396 14724 12430
rect 14539 12391 14724 12396
rect 14539 12357 14609 12391
rect 14643 12358 14724 12391
rect 14539 12324 14614 12357
rect 14648 12324 14724 12358
rect 14539 12323 14724 12324
rect 14539 12289 14609 12323
rect 14643 12289 14724 12323
rect 14539 12286 14724 12289
rect 14539 12255 14614 12286
rect 14539 12221 14609 12255
rect 14648 12252 14724 12286
rect 14643 12221 14724 12252
rect 14539 12214 14724 12221
rect 14539 12187 14614 12214
rect 14539 12153 14609 12187
rect 14648 12180 14724 12214
rect 14643 12153 14724 12180
rect 14539 12142 14724 12153
rect 14539 12119 14614 12142
rect 14539 12085 14609 12119
rect 14648 12108 14724 12142
rect 14643 12085 14724 12108
rect 14539 12070 14724 12085
rect 14539 12051 14614 12070
rect 14539 12017 14609 12051
rect 14648 12036 14724 12070
rect 14643 12017 14724 12036
rect 14539 11998 14724 12017
rect 14539 11983 14614 11998
rect 14539 11949 14609 11983
rect 14648 11964 14724 11998
rect 14643 11949 14724 11964
rect 14539 11926 14724 11949
rect 14539 11915 14614 11926
rect 14539 11881 14609 11915
rect 14648 11892 14724 11926
rect 14643 11881 14724 11892
rect 14539 11854 14724 11881
rect 14539 11847 14614 11854
rect 14539 11813 14609 11847
rect 14648 11820 14724 11854
rect 14643 11813 14724 11820
rect 14539 11782 14724 11813
rect 14539 11779 14614 11782
rect 14539 11745 14609 11779
rect 14648 11748 14724 11782
rect 14643 11745 14724 11748
rect 14539 11711 14724 11745
rect 14539 11677 14609 11711
rect 14643 11710 14724 11711
rect 14539 11676 14614 11677
rect 14648 11676 14724 11710
rect 14539 11643 14724 11676
rect 14539 11609 14609 11643
rect 14643 11638 14724 11643
rect 14539 11604 14614 11609
rect 14648 11604 14724 11638
rect 14539 11575 14724 11604
rect 14539 11541 14609 11575
rect 14643 11566 14724 11575
rect 14539 11532 14614 11541
rect 14648 11532 14724 11566
rect 14539 11507 14724 11532
rect 14539 11473 14609 11507
rect 14643 11494 14724 11507
rect 14539 11460 14614 11473
rect 14648 11460 14724 11494
rect 14539 11439 14724 11460
rect 14539 11405 14609 11439
rect 14643 11422 14724 11439
rect 14539 11388 14614 11405
rect 14648 11388 14724 11422
rect 14539 11371 14724 11388
rect 14539 11337 14609 11371
rect 14643 11350 14724 11371
rect 14539 11316 14614 11337
rect 14648 11316 14724 11350
rect 14539 11303 14724 11316
rect 14539 11269 14609 11303
rect 14643 11278 14724 11303
rect 14539 11244 14614 11269
rect 14648 11244 14724 11278
rect 14539 11235 14724 11244
rect 14539 11201 14609 11235
rect 14643 11206 14724 11235
rect 14539 11172 14614 11201
rect 14648 11172 14724 11206
rect 14539 11167 14724 11172
rect 14539 11133 14609 11167
rect 14643 11134 14724 11167
rect 14539 11100 14614 11133
rect 14648 11100 14724 11134
rect 14539 11099 14724 11100
rect 14539 11065 14609 11099
rect 14643 11065 14724 11099
rect 14539 11062 14724 11065
rect 14539 11031 14614 11062
rect 14539 10997 14609 11031
rect 14648 11028 14724 11062
rect 14643 10997 14724 11028
rect 14539 10990 14724 10997
rect 14539 10963 14614 10990
rect 14539 10929 14609 10963
rect 14648 10956 14724 10990
rect 14643 10929 14724 10956
rect 14539 10918 14724 10929
rect 14539 10895 14614 10918
rect 14539 10861 14609 10895
rect 14648 10884 14724 10918
rect 14643 10861 14724 10884
rect 14539 10846 14724 10861
rect 14539 10827 14614 10846
rect 14539 10793 14609 10827
rect 14648 10812 14724 10846
rect 14643 10793 14724 10812
rect 14539 10774 14724 10793
rect 14539 10759 14614 10774
rect 14539 10725 14609 10759
rect 14648 10740 14724 10774
rect 14643 10725 14724 10740
rect 14539 10702 14724 10725
rect 14539 10691 14614 10702
rect 14539 10657 14609 10691
rect 14648 10668 14724 10702
rect 14643 10657 14724 10668
rect 14539 10630 14724 10657
rect 14539 10623 14614 10630
rect 14539 10589 14609 10623
rect 14648 10596 14724 10630
rect 14643 10589 14724 10596
rect 14539 10558 14724 10589
rect 14539 10555 14614 10558
rect 14539 10521 14609 10555
rect 14648 10524 14724 10558
rect 14643 10521 14724 10524
rect 14539 10487 14724 10521
rect 14539 10453 14609 10487
rect 14643 10486 14724 10487
rect 14539 10452 14614 10453
rect 14648 10452 14724 10486
rect 14539 10419 14724 10452
rect 14539 10385 14609 10419
rect 14643 10414 14724 10419
rect 14539 10380 14614 10385
rect 14648 10380 14724 10414
rect 14539 10351 14724 10380
rect 14539 10317 14609 10351
rect 14643 10342 14724 10351
rect 14539 10308 14614 10317
rect 14648 10308 14724 10342
rect 14539 10283 14724 10308
rect 14539 10249 14609 10283
rect 14643 10270 14724 10283
rect 14539 10236 14614 10249
rect 14648 10236 14724 10270
rect 14539 10215 14724 10236
rect 14539 10181 14609 10215
rect 14643 10198 14724 10215
rect 14539 10164 14614 10181
rect 14648 10164 14724 10198
rect 14539 10147 14724 10164
rect 14539 10113 14609 10147
rect 14643 10126 14724 10147
rect 14539 10092 14614 10113
rect 14648 10092 14724 10126
rect 14539 10079 14724 10092
rect 14539 10045 14609 10079
rect 14643 10054 14724 10079
rect 14539 10020 14614 10045
rect 14648 10020 14724 10054
rect 14539 10011 14724 10020
rect 14539 9977 14609 10011
rect 14643 9982 14724 10011
rect 14539 9948 14614 9977
rect 14648 9948 14724 9982
rect 14539 9943 14724 9948
rect 14539 9909 14609 9943
rect 14643 9910 14724 9943
rect 14539 9876 14614 9909
rect 14648 9876 14724 9910
rect 14539 9875 14724 9876
rect 14539 9841 14609 9875
rect 14643 9841 14724 9875
rect 14539 9838 14724 9841
rect 14539 9807 14614 9838
rect 14539 9773 14609 9807
rect 14648 9804 14724 9838
rect 14643 9773 14724 9804
rect 14539 9766 14724 9773
rect 14539 9739 14614 9766
rect 910 9710 2070 9711
rect 12882 9710 14070 9711
rect 245 9663 320 9697
rect 354 9679 430 9697
rect 245 9645 322 9663
rect 356 9645 430 9679
rect 245 9611 430 9645
rect 245 9577 322 9611
rect 356 9577 430 9611
rect 245 9528 430 9577
rect 14539 9705 14609 9739
rect 14648 9732 14724 9766
rect 14643 9705 14724 9732
rect 14539 9694 14724 9705
rect 14539 9671 14614 9694
rect 14539 9637 14609 9671
rect 14648 9660 14724 9694
rect 14643 9637 14724 9660
rect 14539 9603 14724 9637
rect 14539 9569 14609 9603
rect 14643 9569 14724 9603
rect 14539 9528 14724 9569
rect 245 9454 14724 9528
rect 245 9452 510 9454
rect 245 9418 320 9452
rect 354 9420 510 9452
rect 544 9420 578 9454
rect 612 9452 646 9454
rect 644 9420 646 9452
rect 680 9420 714 9454
rect 748 9420 782 9454
rect 816 9420 850 9454
rect 884 9420 918 9454
rect 952 9420 986 9454
rect 1020 9420 1054 9454
rect 1088 9420 1122 9454
rect 1156 9420 1190 9454
rect 1224 9420 1258 9454
rect 1292 9420 1326 9454
rect 1360 9420 1394 9454
rect 1428 9420 1462 9454
rect 1496 9420 1530 9454
rect 1564 9420 1598 9454
rect 1632 9420 1666 9454
rect 1700 9420 1734 9454
rect 1768 9420 1802 9454
rect 1836 9420 1870 9454
rect 1904 9420 1938 9454
rect 1972 9420 2006 9454
rect 2040 9420 2074 9454
rect 2108 9420 2142 9454
rect 2176 9420 2210 9454
rect 2244 9420 2278 9454
rect 2312 9452 2346 9454
rect 2345 9420 2346 9452
rect 2380 9452 2414 9454
rect 2448 9452 2482 9454
rect 2516 9452 2550 9454
rect 2584 9452 2618 9454
rect 2652 9452 2686 9454
rect 2720 9452 2754 9454
rect 2788 9452 2822 9454
rect 2856 9452 2890 9454
rect 2380 9420 2383 9452
rect 2448 9420 2455 9452
rect 2516 9420 2527 9452
rect 2584 9420 2599 9452
rect 2652 9420 2671 9452
rect 2720 9420 2743 9452
rect 2788 9420 2815 9452
rect 2856 9420 2887 9452
rect 2924 9420 2958 9454
rect 2992 9452 3026 9454
rect 3060 9452 3094 9454
rect 3128 9452 3162 9454
rect 3196 9452 3230 9454
rect 3264 9452 3298 9454
rect 3332 9452 3366 9454
rect 3400 9452 3434 9454
rect 3468 9452 3502 9454
rect 3536 9452 3570 9454
rect 2993 9420 3026 9452
rect 3065 9420 3094 9452
rect 3137 9420 3162 9452
rect 3209 9420 3230 9452
rect 3281 9420 3298 9452
rect 3353 9420 3366 9452
rect 3425 9420 3434 9452
rect 3497 9420 3502 9452
rect 3569 9420 3570 9452
rect 3604 9452 3638 9454
rect 3672 9452 3706 9454
rect 3740 9452 3774 9454
rect 3808 9452 3842 9454
rect 3876 9452 3910 9454
rect 3944 9452 3978 9454
rect 4012 9452 4046 9454
rect 4080 9452 4114 9454
rect 3604 9420 3607 9452
rect 3672 9420 3679 9452
rect 3740 9420 3751 9452
rect 3808 9420 3823 9452
rect 3876 9420 3895 9452
rect 3944 9420 3967 9452
rect 4012 9420 4039 9452
rect 4080 9420 4111 9452
rect 4148 9420 4182 9454
rect 4216 9452 4250 9454
rect 4284 9452 4318 9454
rect 4352 9452 4386 9454
rect 4420 9452 4454 9454
rect 4488 9452 4522 9454
rect 4556 9452 4590 9454
rect 4624 9452 4658 9454
rect 4692 9452 4726 9454
rect 4760 9452 4794 9454
rect 4217 9420 4250 9452
rect 4289 9420 4318 9452
rect 4361 9420 4386 9452
rect 4433 9420 4454 9452
rect 4505 9420 4522 9452
rect 4577 9420 4590 9452
rect 4649 9420 4658 9452
rect 4721 9420 4726 9452
rect 4793 9420 4794 9452
rect 4828 9452 4862 9454
rect 4896 9452 4930 9454
rect 4964 9452 4998 9454
rect 5032 9452 5066 9454
rect 5100 9452 5134 9454
rect 5168 9452 5202 9454
rect 5236 9452 5270 9454
rect 5304 9452 5338 9454
rect 4828 9420 4831 9452
rect 4896 9420 4903 9452
rect 4964 9420 4975 9452
rect 5032 9420 5047 9452
rect 5100 9420 5119 9452
rect 5168 9420 5191 9452
rect 5236 9420 5263 9452
rect 5304 9420 5335 9452
rect 5372 9420 5406 9454
rect 5440 9452 5474 9454
rect 5508 9452 5542 9454
rect 5576 9452 5610 9454
rect 5644 9452 5678 9454
rect 5712 9452 5746 9454
rect 5780 9452 5814 9454
rect 5848 9452 5882 9454
rect 5916 9452 5950 9454
rect 5984 9452 6018 9454
rect 5441 9420 5474 9452
rect 5513 9420 5542 9452
rect 5585 9420 5610 9452
rect 5657 9420 5678 9452
rect 5729 9420 5746 9452
rect 5801 9420 5814 9452
rect 5873 9420 5882 9452
rect 5945 9420 5950 9452
rect 6017 9420 6018 9452
rect 6052 9452 6086 9454
rect 6120 9452 6154 9454
rect 6188 9452 6222 9454
rect 6256 9452 6290 9454
rect 6324 9452 6358 9454
rect 6392 9452 6426 9454
rect 6460 9452 6494 9454
rect 6528 9452 6562 9454
rect 6052 9420 6055 9452
rect 6120 9420 6127 9452
rect 6188 9420 6199 9452
rect 6256 9420 6271 9452
rect 6324 9420 6343 9452
rect 6392 9420 6415 9452
rect 6460 9420 6487 9452
rect 6528 9420 6559 9452
rect 6596 9420 6630 9454
rect 6664 9452 6698 9454
rect 6732 9452 6766 9454
rect 6800 9452 6834 9454
rect 6868 9452 6902 9454
rect 6936 9452 6970 9454
rect 7004 9452 7038 9454
rect 7072 9452 7106 9454
rect 7140 9452 7174 9454
rect 7208 9452 7242 9454
rect 6665 9420 6698 9452
rect 6737 9420 6766 9452
rect 6809 9420 6834 9452
rect 6881 9420 6902 9452
rect 6953 9420 6970 9452
rect 7025 9420 7038 9452
rect 7097 9420 7106 9452
rect 7169 9420 7174 9452
rect 7241 9420 7242 9452
rect 7276 9452 7310 9454
rect 7344 9452 7378 9454
rect 7412 9452 7446 9454
rect 7480 9452 7514 9454
rect 7548 9452 7582 9454
rect 7616 9452 7650 9454
rect 7684 9452 7718 9454
rect 7752 9452 7786 9454
rect 7276 9420 7279 9452
rect 7344 9420 7351 9452
rect 7412 9420 7423 9452
rect 7480 9420 7495 9452
rect 7548 9420 7567 9452
rect 7616 9420 7639 9452
rect 7684 9420 7711 9452
rect 7752 9420 7783 9452
rect 7820 9420 7854 9454
rect 7888 9452 7922 9454
rect 7956 9452 7990 9454
rect 8024 9452 8058 9454
rect 8092 9452 8126 9454
rect 8160 9452 8194 9454
rect 8228 9452 8262 9454
rect 8296 9452 8330 9454
rect 8364 9452 8398 9454
rect 8432 9452 8466 9454
rect 7889 9420 7922 9452
rect 7961 9420 7990 9452
rect 8033 9420 8058 9452
rect 8105 9420 8126 9452
rect 8177 9420 8194 9452
rect 8249 9420 8262 9452
rect 8321 9420 8330 9452
rect 8393 9420 8398 9452
rect 8465 9420 8466 9452
rect 8500 9452 8534 9454
rect 8568 9452 8602 9454
rect 8636 9452 8670 9454
rect 8704 9452 8738 9454
rect 8772 9452 8806 9454
rect 8840 9452 8874 9454
rect 8908 9452 8942 9454
rect 8976 9452 9010 9454
rect 8500 9420 8503 9452
rect 8568 9420 8575 9452
rect 8636 9420 8647 9452
rect 8704 9420 8719 9452
rect 8772 9420 8791 9452
rect 8840 9420 8863 9452
rect 8908 9420 8935 9452
rect 8976 9420 9007 9452
rect 9044 9420 9078 9454
rect 9112 9452 9146 9454
rect 9180 9452 9214 9454
rect 9248 9452 9282 9454
rect 9316 9452 9350 9454
rect 9384 9452 9418 9454
rect 9452 9452 9486 9454
rect 9520 9452 9554 9454
rect 9588 9452 9622 9454
rect 9656 9452 9690 9454
rect 9113 9420 9146 9452
rect 9185 9420 9214 9452
rect 9257 9420 9282 9452
rect 9329 9420 9350 9452
rect 9401 9420 9418 9452
rect 9473 9420 9486 9452
rect 9545 9420 9554 9452
rect 9617 9420 9622 9452
rect 9689 9420 9690 9452
rect 9724 9452 9758 9454
rect 9792 9452 9826 9454
rect 9860 9452 9894 9454
rect 9928 9452 9962 9454
rect 9996 9452 10030 9454
rect 10064 9452 10098 9454
rect 10132 9452 10166 9454
rect 10200 9452 10234 9454
rect 9724 9420 9727 9452
rect 9792 9420 9799 9452
rect 9860 9420 9871 9452
rect 9928 9420 9943 9452
rect 9996 9420 10015 9452
rect 10064 9420 10087 9452
rect 10132 9420 10159 9452
rect 10200 9420 10231 9452
rect 10268 9420 10302 9454
rect 10336 9452 10370 9454
rect 10404 9452 10438 9454
rect 10472 9452 10506 9454
rect 10540 9452 10574 9454
rect 10608 9452 10642 9454
rect 10676 9452 10710 9454
rect 10744 9452 10778 9454
rect 10812 9452 10846 9454
rect 10880 9452 10914 9454
rect 10337 9420 10370 9452
rect 10409 9420 10438 9452
rect 10481 9420 10506 9452
rect 10553 9420 10574 9452
rect 10625 9420 10642 9452
rect 10697 9420 10710 9452
rect 10769 9420 10778 9452
rect 10841 9420 10846 9452
rect 10913 9420 10914 9452
rect 10948 9452 10982 9454
rect 11016 9452 11050 9454
rect 11084 9452 11118 9454
rect 11152 9452 11186 9454
rect 11220 9452 11254 9454
rect 11288 9452 11322 9454
rect 11356 9452 11390 9454
rect 11424 9452 11458 9454
rect 10948 9420 10951 9452
rect 11016 9420 11023 9452
rect 11084 9420 11095 9452
rect 11152 9420 11167 9452
rect 11220 9420 11239 9452
rect 11288 9420 11311 9452
rect 11356 9420 11383 9452
rect 11424 9420 11455 9452
rect 11492 9420 11526 9454
rect 11560 9452 11594 9454
rect 11628 9452 11662 9454
rect 11696 9452 11730 9454
rect 11764 9452 11798 9454
rect 11832 9452 11866 9454
rect 11900 9452 11934 9454
rect 11968 9452 12002 9454
rect 12036 9452 12070 9454
rect 12104 9452 12138 9454
rect 11561 9420 11594 9452
rect 11633 9420 11662 9452
rect 11705 9420 11730 9452
rect 11777 9420 11798 9452
rect 11849 9420 11866 9452
rect 11921 9420 11934 9452
rect 11993 9420 12002 9452
rect 12065 9420 12070 9452
rect 12137 9420 12138 9452
rect 12172 9452 12206 9454
rect 12240 9452 12274 9454
rect 12308 9452 12342 9454
rect 12376 9452 12410 9454
rect 12444 9452 12478 9454
rect 12512 9452 12546 9454
rect 12580 9452 12614 9454
rect 12172 9420 12175 9452
rect 12240 9420 12247 9452
rect 12308 9420 12319 9452
rect 12376 9420 12391 9452
rect 12444 9420 12463 9452
rect 12512 9420 12535 9452
rect 12580 9420 12607 9452
rect 12648 9420 12682 9454
rect 12716 9420 12750 9454
rect 12784 9420 12818 9454
rect 12852 9420 12886 9454
rect 12920 9420 12954 9454
rect 12988 9420 13022 9454
rect 13056 9420 13090 9454
rect 13124 9420 13158 9454
rect 13192 9420 13226 9454
rect 13260 9420 13294 9454
rect 13328 9420 13362 9454
rect 13396 9420 13430 9454
rect 13464 9420 13498 9454
rect 13532 9420 13566 9454
rect 13600 9420 13634 9454
rect 13668 9420 13702 9454
rect 13736 9420 13770 9454
rect 13804 9420 13838 9454
rect 13872 9420 13906 9454
rect 13940 9420 13974 9454
rect 14008 9420 14042 9454
rect 14076 9420 14110 9454
rect 14144 9420 14178 9454
rect 14212 9420 14246 9454
rect 14280 9420 14314 9454
rect 14348 9420 14382 9454
rect 14416 9420 14450 9454
rect 14484 9452 14724 9454
rect 14484 9420 14614 9452
rect 354 9418 610 9420
rect 644 9418 2311 9420
rect 2345 9418 2383 9420
rect 2417 9418 2455 9420
rect 2489 9418 2527 9420
rect 2561 9418 2599 9420
rect 2633 9418 2671 9420
rect 2705 9418 2743 9420
rect 2777 9418 2815 9420
rect 2849 9418 2887 9420
rect 2921 9418 2959 9420
rect 2993 9418 3031 9420
rect 3065 9418 3103 9420
rect 3137 9418 3175 9420
rect 3209 9418 3247 9420
rect 3281 9418 3319 9420
rect 3353 9418 3391 9420
rect 3425 9418 3463 9420
rect 3497 9418 3535 9420
rect 3569 9418 3607 9420
rect 3641 9418 3679 9420
rect 3713 9418 3751 9420
rect 3785 9418 3823 9420
rect 3857 9418 3895 9420
rect 3929 9418 3967 9420
rect 4001 9418 4039 9420
rect 4073 9418 4111 9420
rect 4145 9418 4183 9420
rect 4217 9418 4255 9420
rect 4289 9418 4327 9420
rect 4361 9418 4399 9420
rect 4433 9418 4471 9420
rect 4505 9418 4543 9420
rect 4577 9418 4615 9420
rect 4649 9418 4687 9420
rect 4721 9418 4759 9420
rect 4793 9418 4831 9420
rect 4865 9418 4903 9420
rect 4937 9418 4975 9420
rect 5009 9418 5047 9420
rect 5081 9418 5119 9420
rect 5153 9418 5191 9420
rect 5225 9418 5263 9420
rect 5297 9418 5335 9420
rect 5369 9418 5407 9420
rect 5441 9418 5479 9420
rect 5513 9418 5551 9420
rect 5585 9418 5623 9420
rect 5657 9418 5695 9420
rect 5729 9418 5767 9420
rect 5801 9418 5839 9420
rect 5873 9418 5911 9420
rect 5945 9418 5983 9420
rect 6017 9418 6055 9420
rect 6089 9418 6127 9420
rect 6161 9418 6199 9420
rect 6233 9418 6271 9420
rect 6305 9418 6343 9420
rect 6377 9418 6415 9420
rect 6449 9418 6487 9420
rect 6521 9418 6559 9420
rect 6593 9418 6631 9420
rect 6665 9418 6703 9420
rect 6737 9418 6775 9420
rect 6809 9418 6847 9420
rect 6881 9418 6919 9420
rect 6953 9418 6991 9420
rect 7025 9418 7063 9420
rect 7097 9418 7135 9420
rect 7169 9418 7207 9420
rect 7241 9418 7279 9420
rect 7313 9418 7351 9420
rect 7385 9418 7423 9420
rect 7457 9418 7495 9420
rect 7529 9418 7567 9420
rect 7601 9418 7639 9420
rect 7673 9418 7711 9420
rect 7745 9418 7783 9420
rect 7817 9418 7855 9420
rect 7889 9418 7927 9420
rect 7961 9418 7999 9420
rect 8033 9418 8071 9420
rect 8105 9418 8143 9420
rect 8177 9418 8215 9420
rect 8249 9418 8287 9420
rect 8321 9418 8359 9420
rect 8393 9418 8431 9420
rect 8465 9418 8503 9420
rect 8537 9418 8575 9420
rect 8609 9418 8647 9420
rect 8681 9418 8719 9420
rect 8753 9418 8791 9420
rect 8825 9418 8863 9420
rect 8897 9418 8935 9420
rect 8969 9418 9007 9420
rect 9041 9418 9079 9420
rect 9113 9418 9151 9420
rect 9185 9418 9223 9420
rect 9257 9418 9295 9420
rect 9329 9418 9367 9420
rect 9401 9418 9439 9420
rect 9473 9418 9511 9420
rect 9545 9418 9583 9420
rect 9617 9418 9655 9420
rect 9689 9418 9727 9420
rect 9761 9418 9799 9420
rect 9833 9418 9871 9420
rect 9905 9418 9943 9420
rect 9977 9418 10015 9420
rect 10049 9418 10087 9420
rect 10121 9418 10159 9420
rect 10193 9418 10231 9420
rect 10265 9418 10303 9420
rect 10337 9418 10375 9420
rect 10409 9418 10447 9420
rect 10481 9418 10519 9420
rect 10553 9418 10591 9420
rect 10625 9418 10663 9420
rect 10697 9418 10735 9420
rect 10769 9418 10807 9420
rect 10841 9418 10879 9420
rect 10913 9418 10951 9420
rect 10985 9418 11023 9420
rect 11057 9418 11095 9420
rect 11129 9418 11167 9420
rect 11201 9418 11239 9420
rect 11273 9418 11311 9420
rect 11345 9418 11383 9420
rect 11417 9418 11455 9420
rect 11489 9418 11527 9420
rect 11561 9418 11599 9420
rect 11633 9418 11671 9420
rect 11705 9418 11743 9420
rect 11777 9418 11815 9420
rect 11849 9418 11887 9420
rect 11921 9418 11959 9420
rect 11993 9418 12031 9420
rect 12065 9418 12103 9420
rect 12137 9418 12175 9420
rect 12209 9418 12247 9420
rect 12281 9418 12319 9420
rect 12353 9418 12391 9420
rect 12425 9418 12463 9420
rect 12497 9418 12535 9420
rect 12569 9418 12607 9420
rect 12641 9418 14314 9420
rect 14348 9418 14614 9420
rect 14648 9418 14724 9452
rect 245 9343 14724 9418
<< viali >>
rect 320 36500 354 36534
rect 14614 36499 14648 36533
rect 556 36465 560 36498
rect 560 36465 590 36498
rect 628 36465 662 36498
rect 700 36465 730 36498
rect 730 36465 734 36498
rect 772 36465 798 36498
rect 798 36465 806 36498
rect 844 36465 866 36498
rect 866 36465 878 36498
rect 916 36465 934 36498
rect 934 36465 950 36498
rect 988 36465 1002 36498
rect 1002 36465 1022 36498
rect 1060 36465 1070 36498
rect 1070 36465 1094 36498
rect 1132 36465 1138 36498
rect 1138 36465 1166 36498
rect 1204 36465 1206 36498
rect 1206 36465 1238 36498
rect 1276 36465 1308 36498
rect 1308 36465 1310 36498
rect 1348 36465 1376 36498
rect 1376 36465 1382 36498
rect 1420 36465 1444 36498
rect 1444 36465 1454 36498
rect 1492 36465 1512 36498
rect 1512 36465 1526 36498
rect 1564 36465 1580 36498
rect 1580 36465 1598 36498
rect 1636 36465 1648 36498
rect 1648 36465 1670 36498
rect 1708 36465 1716 36498
rect 1716 36465 1742 36498
rect 1780 36465 1784 36498
rect 1784 36465 1814 36498
rect 1852 36465 1886 36498
rect 1924 36465 1954 36498
rect 1954 36465 1958 36498
rect 1996 36465 2022 36498
rect 2022 36465 2030 36498
rect 2068 36465 2090 36498
rect 2090 36465 2102 36498
rect 2140 36465 2158 36498
rect 2158 36465 2174 36498
rect 2212 36465 2226 36498
rect 2226 36465 2246 36498
rect 2284 36465 2294 36498
rect 2294 36465 2318 36498
rect 2356 36465 2362 36498
rect 2362 36465 2390 36498
rect 2428 36465 2430 36498
rect 2430 36465 2462 36498
rect 2500 36465 2532 36498
rect 2532 36465 2534 36498
rect 2572 36465 2600 36498
rect 2600 36465 2606 36498
rect 2644 36465 2668 36498
rect 2668 36465 2678 36498
rect 2716 36465 2736 36498
rect 2736 36465 2750 36498
rect 2788 36465 2804 36498
rect 2804 36465 2822 36498
rect 2860 36465 2872 36498
rect 2872 36465 2894 36498
rect 2932 36465 2940 36498
rect 2940 36465 2966 36498
rect 3004 36465 3008 36498
rect 3008 36465 3038 36498
rect 3076 36465 3110 36498
rect 3148 36465 3178 36498
rect 3178 36465 3182 36498
rect 3220 36465 3246 36498
rect 3246 36465 3254 36498
rect 3292 36465 3314 36498
rect 3314 36465 3326 36498
rect 3364 36465 3382 36498
rect 3382 36465 3398 36498
rect 3436 36465 3450 36498
rect 3450 36465 3470 36498
rect 3508 36465 3518 36498
rect 3518 36465 3542 36498
rect 3580 36465 3586 36498
rect 3586 36465 3614 36498
rect 3652 36465 3654 36498
rect 3654 36465 3686 36498
rect 3724 36465 3756 36498
rect 3756 36465 3758 36498
rect 3796 36465 3824 36498
rect 3824 36465 3830 36498
rect 3868 36465 3892 36498
rect 3892 36465 3902 36498
rect 3940 36465 3960 36498
rect 3960 36465 3974 36498
rect 4012 36465 4028 36498
rect 4028 36465 4046 36498
rect 4084 36465 4096 36498
rect 4096 36465 4118 36498
rect 4156 36465 4164 36498
rect 4164 36465 4190 36498
rect 4228 36465 4232 36498
rect 4232 36465 4262 36498
rect 4300 36465 4334 36498
rect 4372 36465 4402 36498
rect 4402 36465 4406 36498
rect 4444 36465 4470 36498
rect 4470 36465 4478 36498
rect 4516 36465 4538 36498
rect 4538 36465 4550 36498
rect 4588 36465 4606 36498
rect 4606 36465 4622 36498
rect 4660 36465 4674 36498
rect 4674 36465 4694 36498
rect 4732 36465 4742 36498
rect 4742 36465 4766 36498
rect 4804 36465 4810 36498
rect 4810 36465 4838 36498
rect 4876 36465 4878 36498
rect 4878 36465 4910 36498
rect 4948 36465 4980 36498
rect 4980 36465 4982 36498
rect 5020 36465 5048 36498
rect 5048 36465 5054 36498
rect 5092 36465 5116 36498
rect 5116 36465 5126 36498
rect 5164 36465 5184 36498
rect 5184 36465 5198 36498
rect 5236 36465 5252 36498
rect 5252 36465 5270 36498
rect 5308 36465 5320 36498
rect 5320 36465 5342 36498
rect 5380 36465 5388 36498
rect 5388 36465 5414 36498
rect 5452 36465 5456 36498
rect 5456 36465 5486 36498
rect 5524 36465 5558 36498
rect 5596 36465 5626 36498
rect 5626 36465 5630 36498
rect 5668 36465 5694 36498
rect 5694 36465 5702 36498
rect 5740 36465 5762 36498
rect 5762 36465 5774 36498
rect 5812 36465 5830 36498
rect 5830 36465 5846 36498
rect 5884 36465 5898 36498
rect 5898 36465 5918 36498
rect 5956 36465 5966 36498
rect 5966 36465 5990 36498
rect 6028 36465 6034 36498
rect 6034 36465 6062 36498
rect 6100 36465 6102 36498
rect 6102 36465 6134 36498
rect 6172 36465 6204 36498
rect 6204 36465 6206 36498
rect 6244 36465 6272 36498
rect 6272 36465 6278 36498
rect 6316 36465 6340 36498
rect 6340 36465 6350 36498
rect 6388 36465 6408 36498
rect 6408 36465 6422 36498
rect 6460 36465 6476 36498
rect 6476 36465 6494 36498
rect 6532 36465 6544 36498
rect 6544 36465 6566 36498
rect 6604 36465 6612 36498
rect 6612 36465 6638 36498
rect 6676 36465 6680 36498
rect 6680 36465 6710 36498
rect 6748 36465 6782 36498
rect 6820 36465 6850 36498
rect 6850 36465 6854 36498
rect 6892 36465 6918 36498
rect 6918 36465 6926 36498
rect 6964 36465 6986 36498
rect 6986 36465 6998 36498
rect 7036 36465 7054 36498
rect 7054 36465 7070 36498
rect 7108 36465 7122 36498
rect 7122 36465 7142 36498
rect 7180 36465 7190 36498
rect 7190 36465 7214 36498
rect 7252 36465 7258 36498
rect 7258 36465 7286 36498
rect 7324 36465 7326 36498
rect 7326 36465 7358 36498
rect 7396 36465 7428 36498
rect 7428 36465 7430 36498
rect 7468 36465 7496 36498
rect 7496 36465 7502 36498
rect 7540 36465 7564 36498
rect 7564 36465 7574 36498
rect 7612 36465 7632 36498
rect 7632 36465 7646 36498
rect 7684 36465 7700 36498
rect 7700 36465 7718 36498
rect 7756 36465 7768 36498
rect 7768 36465 7790 36498
rect 7828 36465 7836 36498
rect 7836 36465 7862 36498
rect 7900 36465 7904 36498
rect 7904 36465 7934 36498
rect 7972 36465 8006 36498
rect 8044 36465 8074 36498
rect 8074 36465 8078 36498
rect 8116 36465 8142 36498
rect 8142 36465 8150 36498
rect 8188 36465 8210 36498
rect 8210 36465 8222 36498
rect 8260 36465 8278 36498
rect 8278 36465 8294 36498
rect 8332 36465 8346 36498
rect 8346 36465 8366 36498
rect 8404 36465 8414 36498
rect 8414 36465 8438 36498
rect 8476 36465 8482 36498
rect 8482 36465 8510 36498
rect 8548 36465 8550 36498
rect 8550 36465 8582 36498
rect 8620 36465 8652 36498
rect 8652 36465 8654 36498
rect 8692 36465 8720 36498
rect 8720 36465 8726 36498
rect 8764 36465 8788 36498
rect 8788 36465 8798 36498
rect 8836 36465 8856 36498
rect 8856 36465 8870 36498
rect 8908 36465 8924 36498
rect 8924 36465 8942 36498
rect 8980 36465 8992 36498
rect 8992 36465 9014 36498
rect 9052 36465 9060 36498
rect 9060 36465 9086 36498
rect 9124 36465 9128 36498
rect 9128 36465 9158 36498
rect 9196 36465 9230 36498
rect 9268 36465 9298 36498
rect 9298 36465 9302 36498
rect 9340 36465 9366 36498
rect 9366 36465 9374 36498
rect 9412 36465 9434 36498
rect 9434 36465 9446 36498
rect 9484 36465 9502 36498
rect 9502 36465 9518 36498
rect 9556 36465 9570 36498
rect 9570 36465 9590 36498
rect 9628 36465 9638 36498
rect 9638 36465 9662 36498
rect 9700 36465 9706 36498
rect 9706 36465 9734 36498
rect 9772 36465 9774 36498
rect 9774 36465 9806 36498
rect 9844 36465 9876 36498
rect 9876 36465 9878 36498
rect 9916 36465 9944 36498
rect 9944 36465 9950 36498
rect 9988 36465 10012 36498
rect 10012 36465 10022 36498
rect 10060 36465 10080 36498
rect 10080 36465 10094 36498
rect 10132 36465 10148 36498
rect 10148 36465 10166 36498
rect 10204 36465 10216 36498
rect 10216 36465 10238 36498
rect 10276 36465 10284 36498
rect 10284 36465 10310 36498
rect 10348 36465 10352 36498
rect 10352 36465 10382 36498
rect 10420 36465 10454 36498
rect 10492 36465 10522 36498
rect 10522 36465 10526 36498
rect 10564 36465 10590 36498
rect 10590 36465 10598 36498
rect 10636 36465 10658 36498
rect 10658 36465 10670 36498
rect 10708 36465 10726 36498
rect 10726 36465 10742 36498
rect 10780 36465 10794 36498
rect 10794 36465 10814 36498
rect 10852 36465 10862 36498
rect 10862 36465 10886 36498
rect 10924 36465 10930 36498
rect 10930 36465 10958 36498
rect 10996 36465 10998 36498
rect 10998 36465 11030 36498
rect 11068 36465 11100 36498
rect 11100 36465 11102 36498
rect 11140 36465 11168 36498
rect 11168 36465 11174 36498
rect 11212 36465 11236 36498
rect 11236 36465 11246 36498
rect 11284 36465 11304 36498
rect 11304 36465 11318 36498
rect 11356 36465 11372 36498
rect 11372 36465 11390 36498
rect 11428 36465 11440 36498
rect 11440 36465 11462 36498
rect 11500 36465 11508 36498
rect 11508 36465 11534 36498
rect 11572 36465 11576 36498
rect 11576 36465 11606 36498
rect 11644 36465 11678 36498
rect 11716 36465 11746 36498
rect 11746 36465 11750 36498
rect 11788 36465 11814 36498
rect 11814 36465 11822 36498
rect 11860 36465 11882 36498
rect 11882 36465 11894 36498
rect 11932 36465 11950 36498
rect 11950 36465 11966 36498
rect 12004 36465 12018 36498
rect 12018 36465 12038 36498
rect 12076 36465 12086 36498
rect 12086 36465 12110 36498
rect 12148 36465 12154 36498
rect 12154 36465 12182 36498
rect 12220 36465 12222 36498
rect 12222 36465 12254 36498
rect 12292 36465 12324 36498
rect 12324 36465 12326 36498
rect 12364 36465 12392 36498
rect 12392 36465 12398 36498
rect 12436 36465 12460 36498
rect 12460 36465 12470 36498
rect 12508 36465 12528 36498
rect 12528 36465 12542 36498
rect 12580 36465 12596 36498
rect 12596 36465 12614 36498
rect 12652 36465 12664 36498
rect 12664 36465 12686 36498
rect 12724 36465 12732 36498
rect 12732 36465 12758 36498
rect 12796 36465 12800 36498
rect 12800 36465 12830 36498
rect 12868 36465 12902 36498
rect 12940 36465 12970 36498
rect 12970 36465 12974 36498
rect 13012 36465 13038 36498
rect 13038 36465 13046 36498
rect 13084 36465 13106 36498
rect 13106 36465 13118 36498
rect 13156 36465 13174 36498
rect 13174 36465 13190 36498
rect 13228 36465 13242 36498
rect 13242 36465 13262 36498
rect 13300 36465 13310 36498
rect 13310 36465 13334 36498
rect 13372 36465 13378 36498
rect 13378 36465 13406 36498
rect 13444 36465 13446 36498
rect 13446 36465 13478 36498
rect 13516 36465 13548 36498
rect 13548 36465 13550 36498
rect 13588 36465 13616 36498
rect 13616 36465 13622 36498
rect 13660 36465 13684 36498
rect 13684 36465 13694 36498
rect 13732 36465 13752 36498
rect 13752 36465 13766 36498
rect 13804 36465 13820 36498
rect 13820 36465 13838 36498
rect 13876 36465 13888 36498
rect 13888 36465 13910 36498
rect 13948 36465 13956 36498
rect 13956 36465 13982 36498
rect 14020 36465 14024 36498
rect 14024 36465 14054 36498
rect 14092 36465 14126 36498
rect 14164 36465 14194 36498
rect 14194 36465 14198 36498
rect 14236 36465 14262 36498
rect 14262 36465 14270 36498
rect 14308 36465 14330 36498
rect 14330 36465 14342 36498
rect 14380 36465 14398 36498
rect 14398 36465 14414 36498
rect 556 36464 590 36465
rect 628 36464 662 36465
rect 700 36464 734 36465
rect 772 36464 806 36465
rect 844 36464 878 36465
rect 916 36464 950 36465
rect 988 36464 1022 36465
rect 1060 36464 1094 36465
rect 1132 36464 1166 36465
rect 1204 36464 1238 36465
rect 1276 36464 1310 36465
rect 1348 36464 1382 36465
rect 1420 36464 1454 36465
rect 1492 36464 1526 36465
rect 1564 36464 1598 36465
rect 1636 36464 1670 36465
rect 1708 36464 1742 36465
rect 1780 36464 1814 36465
rect 1852 36464 1886 36465
rect 1924 36464 1958 36465
rect 1996 36464 2030 36465
rect 2068 36464 2102 36465
rect 2140 36464 2174 36465
rect 2212 36464 2246 36465
rect 2284 36464 2318 36465
rect 2356 36464 2390 36465
rect 2428 36464 2462 36465
rect 2500 36464 2534 36465
rect 2572 36464 2606 36465
rect 2644 36464 2678 36465
rect 2716 36464 2750 36465
rect 2788 36464 2822 36465
rect 2860 36464 2894 36465
rect 2932 36464 2966 36465
rect 3004 36464 3038 36465
rect 3076 36464 3110 36465
rect 3148 36464 3182 36465
rect 3220 36464 3254 36465
rect 3292 36464 3326 36465
rect 3364 36464 3398 36465
rect 3436 36464 3470 36465
rect 3508 36464 3542 36465
rect 3580 36464 3614 36465
rect 3652 36464 3686 36465
rect 3724 36464 3758 36465
rect 3796 36464 3830 36465
rect 3868 36464 3902 36465
rect 3940 36464 3974 36465
rect 4012 36464 4046 36465
rect 4084 36464 4118 36465
rect 4156 36464 4190 36465
rect 4228 36464 4262 36465
rect 4300 36464 4334 36465
rect 4372 36464 4406 36465
rect 4444 36464 4478 36465
rect 4516 36464 4550 36465
rect 4588 36464 4622 36465
rect 4660 36464 4694 36465
rect 4732 36464 4766 36465
rect 4804 36464 4838 36465
rect 4876 36464 4910 36465
rect 4948 36464 4982 36465
rect 5020 36464 5054 36465
rect 5092 36464 5126 36465
rect 5164 36464 5198 36465
rect 5236 36464 5270 36465
rect 5308 36464 5342 36465
rect 5380 36464 5414 36465
rect 5452 36464 5486 36465
rect 5524 36464 5558 36465
rect 5596 36464 5630 36465
rect 5668 36464 5702 36465
rect 5740 36464 5774 36465
rect 5812 36464 5846 36465
rect 5884 36464 5918 36465
rect 5956 36464 5990 36465
rect 6028 36464 6062 36465
rect 6100 36464 6134 36465
rect 6172 36464 6206 36465
rect 6244 36464 6278 36465
rect 6316 36464 6350 36465
rect 6388 36464 6422 36465
rect 6460 36464 6494 36465
rect 6532 36464 6566 36465
rect 6604 36464 6638 36465
rect 6676 36464 6710 36465
rect 6748 36464 6782 36465
rect 6820 36464 6854 36465
rect 6892 36464 6926 36465
rect 6964 36464 6998 36465
rect 7036 36464 7070 36465
rect 7108 36464 7142 36465
rect 7180 36464 7214 36465
rect 7252 36464 7286 36465
rect 7324 36464 7358 36465
rect 7396 36464 7430 36465
rect 7468 36464 7502 36465
rect 7540 36464 7574 36465
rect 7612 36464 7646 36465
rect 7684 36464 7718 36465
rect 7756 36464 7790 36465
rect 7828 36464 7862 36465
rect 7900 36464 7934 36465
rect 7972 36464 8006 36465
rect 8044 36464 8078 36465
rect 8116 36464 8150 36465
rect 8188 36464 8222 36465
rect 8260 36464 8294 36465
rect 8332 36464 8366 36465
rect 8404 36464 8438 36465
rect 8476 36464 8510 36465
rect 8548 36464 8582 36465
rect 8620 36464 8654 36465
rect 8692 36464 8726 36465
rect 8764 36464 8798 36465
rect 8836 36464 8870 36465
rect 8908 36464 8942 36465
rect 8980 36464 9014 36465
rect 9052 36464 9086 36465
rect 9124 36464 9158 36465
rect 9196 36464 9230 36465
rect 9268 36464 9302 36465
rect 9340 36464 9374 36465
rect 9412 36464 9446 36465
rect 9484 36464 9518 36465
rect 9556 36464 9590 36465
rect 9628 36464 9662 36465
rect 9700 36464 9734 36465
rect 9772 36464 9806 36465
rect 9844 36464 9878 36465
rect 9916 36464 9950 36465
rect 9988 36464 10022 36465
rect 10060 36464 10094 36465
rect 10132 36464 10166 36465
rect 10204 36464 10238 36465
rect 10276 36464 10310 36465
rect 10348 36464 10382 36465
rect 10420 36464 10454 36465
rect 10492 36464 10526 36465
rect 10564 36464 10598 36465
rect 10636 36464 10670 36465
rect 10708 36464 10742 36465
rect 10780 36464 10814 36465
rect 10852 36464 10886 36465
rect 10924 36464 10958 36465
rect 10996 36464 11030 36465
rect 11068 36464 11102 36465
rect 11140 36464 11174 36465
rect 11212 36464 11246 36465
rect 11284 36464 11318 36465
rect 11356 36464 11390 36465
rect 11428 36464 11462 36465
rect 11500 36464 11534 36465
rect 11572 36464 11606 36465
rect 11644 36464 11678 36465
rect 11716 36464 11750 36465
rect 11788 36464 11822 36465
rect 11860 36464 11894 36465
rect 11932 36464 11966 36465
rect 12004 36464 12038 36465
rect 12076 36464 12110 36465
rect 12148 36464 12182 36465
rect 12220 36464 12254 36465
rect 12292 36464 12326 36465
rect 12364 36464 12398 36465
rect 12436 36464 12470 36465
rect 12508 36464 12542 36465
rect 12580 36464 12614 36465
rect 12652 36464 12686 36465
rect 12724 36464 12758 36465
rect 12796 36464 12830 36465
rect 12868 36464 12902 36465
rect 12940 36464 12974 36465
rect 13012 36464 13046 36465
rect 13084 36464 13118 36465
rect 13156 36464 13190 36465
rect 13228 36464 13262 36465
rect 13300 36464 13334 36465
rect 13372 36464 13406 36465
rect 13444 36464 13478 36465
rect 13516 36464 13550 36465
rect 13588 36464 13622 36465
rect 13660 36464 13694 36465
rect 13732 36464 13766 36465
rect 13804 36464 13838 36465
rect 13876 36464 13910 36465
rect 13948 36464 13982 36465
rect 14020 36464 14054 36465
rect 14092 36464 14126 36465
rect 14164 36464 14198 36465
rect 14236 36464 14270 36465
rect 14308 36464 14342 36465
rect 14380 36464 14414 36465
rect 320 36428 354 36462
rect 14614 36427 14648 36461
rect 320 36233 322 36265
rect 322 36233 354 36265
rect 320 36231 354 36233
rect 14614 36259 14648 36262
rect 14614 36228 14643 36259
rect 14643 36228 14648 36259
rect 320 36165 322 36193
rect 322 36165 354 36193
rect 320 36159 354 36165
rect 320 36097 322 36121
rect 322 36097 354 36121
rect 320 36087 354 36097
rect 320 36029 322 36049
rect 322 36029 354 36049
rect 320 36015 354 36029
rect 320 35961 322 35977
rect 322 35961 354 35977
rect 320 35943 354 35961
rect 320 35893 322 35905
rect 322 35893 354 35905
rect 320 35871 354 35893
rect 320 35825 322 35833
rect 322 35825 354 35833
rect 320 35799 354 35825
rect 320 35757 322 35761
rect 322 35757 354 35761
rect 320 35727 354 35757
rect 320 35655 354 35689
rect 320 35587 354 35617
rect 320 35583 322 35587
rect 322 35583 354 35587
rect 320 35519 354 35545
rect 320 35511 322 35519
rect 322 35511 354 35519
rect 320 35451 354 35473
rect 320 35439 322 35451
rect 322 35439 354 35451
rect 320 35383 354 35401
rect 320 35367 322 35383
rect 322 35367 354 35383
rect 320 35315 354 35329
rect 320 35295 322 35315
rect 322 35295 354 35315
rect 320 35247 354 35257
rect 320 35223 322 35247
rect 322 35223 354 35247
rect 320 35179 354 35185
rect 320 35151 322 35179
rect 322 35151 354 35179
rect 320 35111 354 35113
rect 320 35079 322 35111
rect 322 35079 354 35111
rect 320 35009 322 35041
rect 322 35009 354 35041
rect 320 35007 354 35009
rect 320 34941 322 34969
rect 322 34941 354 34969
rect 320 34935 354 34941
rect 320 34873 322 34897
rect 322 34873 354 34897
rect 320 34863 354 34873
rect 320 34805 322 34825
rect 322 34805 354 34825
rect 320 34791 354 34805
rect 320 34737 322 34753
rect 322 34737 354 34753
rect 320 34719 354 34737
rect 320 34669 322 34681
rect 322 34669 354 34681
rect 320 34647 354 34669
rect 320 34601 322 34609
rect 322 34601 354 34609
rect 320 34575 354 34601
rect 320 34533 322 34537
rect 322 34533 354 34537
rect 320 34503 354 34533
rect 320 34431 354 34465
rect 320 34363 354 34393
rect 320 34359 322 34363
rect 322 34359 354 34363
rect 320 34295 354 34321
rect 320 34287 322 34295
rect 322 34287 354 34295
rect 320 34227 354 34249
rect 320 34215 322 34227
rect 322 34215 354 34227
rect 320 34159 354 34177
rect 320 34143 322 34159
rect 322 34143 354 34159
rect 320 34091 354 34105
rect 320 34071 322 34091
rect 322 34071 354 34091
rect 320 34023 354 34033
rect 320 33999 322 34023
rect 322 33999 354 34023
rect 320 33955 354 33961
rect 320 33927 322 33955
rect 322 33927 354 33955
rect 320 33887 354 33889
rect 320 33855 322 33887
rect 322 33855 354 33887
rect 320 33785 322 33817
rect 322 33785 354 33817
rect 320 33783 354 33785
rect 320 33717 322 33745
rect 322 33717 354 33745
rect 320 33711 354 33717
rect 320 33649 322 33673
rect 322 33649 354 33673
rect 320 33639 354 33649
rect 320 33581 322 33601
rect 322 33581 354 33601
rect 320 33567 354 33581
rect 320 33513 322 33529
rect 322 33513 354 33529
rect 320 33495 354 33513
rect 320 33445 322 33457
rect 322 33445 354 33457
rect 320 33423 354 33445
rect 320 33377 322 33385
rect 322 33377 354 33385
rect 320 33351 354 33377
rect 320 33309 322 33313
rect 322 33309 354 33313
rect 320 33279 354 33309
rect 320 33207 354 33241
rect 320 33139 354 33169
rect 320 33135 322 33139
rect 322 33135 354 33139
rect 320 33071 354 33097
rect 320 33063 322 33071
rect 322 33063 354 33071
rect 320 33003 354 33025
rect 320 32991 322 33003
rect 322 32991 354 33003
rect 320 32935 354 32953
rect 320 32919 322 32935
rect 322 32919 354 32935
rect 320 32867 354 32881
rect 320 32847 322 32867
rect 322 32847 354 32867
rect 320 32799 354 32809
rect 320 32775 322 32799
rect 322 32775 354 32799
rect 320 32731 354 32737
rect 320 32703 322 32731
rect 322 32703 354 32731
rect 320 32663 354 32665
rect 320 32631 322 32663
rect 322 32631 354 32663
rect 320 32561 322 32593
rect 322 32561 354 32593
rect 320 32559 354 32561
rect 320 32493 322 32521
rect 322 32493 354 32521
rect 320 32487 354 32493
rect 320 32425 322 32449
rect 322 32425 354 32449
rect 320 32415 354 32425
rect 320 32357 322 32377
rect 322 32357 354 32377
rect 320 32343 354 32357
rect 320 32289 322 32305
rect 322 32289 354 32305
rect 320 32271 354 32289
rect 320 32221 322 32233
rect 322 32221 354 32233
rect 320 32199 354 32221
rect 320 32153 322 32161
rect 322 32153 354 32161
rect 320 32127 354 32153
rect 320 32085 322 32089
rect 322 32085 354 32089
rect 320 32055 354 32085
rect 320 31983 354 32017
rect 320 31915 354 31945
rect 320 31911 322 31915
rect 322 31911 354 31915
rect 320 31847 354 31873
rect 320 31839 322 31847
rect 322 31839 354 31847
rect 320 31779 354 31801
rect 320 31767 322 31779
rect 322 31767 354 31779
rect 320 31711 354 31729
rect 320 31695 322 31711
rect 322 31695 354 31711
rect 320 31643 354 31657
rect 320 31623 322 31643
rect 322 31623 354 31643
rect 320 31575 354 31585
rect 320 31551 322 31575
rect 322 31551 354 31575
rect 320 31507 354 31513
rect 320 31479 322 31507
rect 322 31479 354 31507
rect 320 31439 354 31441
rect 320 31407 322 31439
rect 322 31407 354 31439
rect 320 31337 322 31369
rect 322 31337 354 31369
rect 320 31335 354 31337
rect 320 31269 322 31297
rect 322 31269 354 31297
rect 320 31263 354 31269
rect 320 31201 322 31225
rect 322 31201 354 31225
rect 320 31191 354 31201
rect 320 31133 322 31153
rect 322 31133 354 31153
rect 320 31119 354 31133
rect 320 31065 322 31081
rect 322 31065 354 31081
rect 320 31047 354 31065
rect 320 30997 322 31009
rect 322 30997 354 31009
rect 320 30975 354 30997
rect 320 30929 322 30937
rect 322 30929 354 30937
rect 320 30903 354 30929
rect 320 30861 322 30865
rect 322 30861 354 30865
rect 320 30831 354 30861
rect 320 30759 354 30793
rect 320 30691 354 30721
rect 320 30687 322 30691
rect 322 30687 354 30691
rect 320 30623 354 30649
rect 320 30615 322 30623
rect 322 30615 354 30623
rect 320 30555 354 30577
rect 320 30543 322 30555
rect 322 30543 354 30555
rect 320 30487 354 30505
rect 320 30471 322 30487
rect 322 30471 354 30487
rect 320 30419 354 30433
rect 320 30399 322 30419
rect 322 30399 354 30419
rect 320 30351 354 30361
rect 320 30327 322 30351
rect 322 30327 354 30351
rect 320 30283 354 30289
rect 320 30255 322 30283
rect 322 30255 354 30283
rect 320 30215 354 30217
rect 320 30183 322 30215
rect 322 30183 354 30215
rect 320 30113 322 30145
rect 322 30113 354 30145
rect 320 30111 354 30113
rect 320 30045 322 30073
rect 322 30045 354 30073
rect 320 30039 354 30045
rect 320 29977 322 30001
rect 322 29977 354 30001
rect 320 29967 354 29977
rect 320 29909 322 29929
rect 322 29909 354 29929
rect 320 29895 354 29909
rect 320 29841 322 29857
rect 322 29841 354 29857
rect 320 29823 354 29841
rect 320 29773 322 29785
rect 322 29773 354 29785
rect 320 29751 354 29773
rect 320 29705 322 29713
rect 322 29705 354 29713
rect 320 29679 354 29705
rect 320 29637 322 29641
rect 322 29637 354 29641
rect 320 29607 354 29637
rect 320 29535 354 29569
rect 320 29467 354 29497
rect 320 29463 322 29467
rect 322 29463 354 29467
rect 320 29399 354 29425
rect 320 29391 322 29399
rect 322 29391 354 29399
rect 320 29331 354 29353
rect 320 29319 322 29331
rect 322 29319 354 29331
rect 320 29263 354 29281
rect 320 29247 322 29263
rect 322 29247 354 29263
rect 320 29195 354 29209
rect 320 29175 322 29195
rect 322 29175 354 29195
rect 320 29127 354 29137
rect 320 29103 322 29127
rect 322 29103 354 29127
rect 320 29059 354 29065
rect 320 29031 322 29059
rect 322 29031 354 29059
rect 320 28991 354 28993
rect 320 28959 322 28991
rect 322 28959 354 28991
rect 320 28889 322 28921
rect 322 28889 354 28921
rect 320 28887 354 28889
rect 320 28821 322 28849
rect 322 28821 354 28849
rect 320 28815 354 28821
rect 320 28753 322 28777
rect 322 28753 354 28777
rect 320 28743 354 28753
rect 320 28685 322 28705
rect 322 28685 354 28705
rect 320 28671 354 28685
rect 320 28617 322 28633
rect 322 28617 354 28633
rect 320 28599 354 28617
rect 320 28549 322 28561
rect 322 28549 354 28561
rect 320 28527 354 28549
rect 320 28481 322 28489
rect 322 28481 354 28489
rect 320 28455 354 28481
rect 320 28413 322 28417
rect 322 28413 354 28417
rect 320 28383 354 28413
rect 320 28311 354 28345
rect 320 28243 354 28273
rect 320 28239 322 28243
rect 322 28239 354 28243
rect 320 28175 354 28201
rect 320 28167 322 28175
rect 322 28167 354 28175
rect 320 28107 354 28129
rect 320 28095 322 28107
rect 322 28095 354 28107
rect 320 28039 354 28057
rect 320 28023 322 28039
rect 322 28023 354 28039
rect 320 27971 354 27985
rect 320 27951 322 27971
rect 322 27951 354 27971
rect 320 27903 354 27913
rect 320 27879 322 27903
rect 322 27879 354 27903
rect 320 27835 354 27841
rect 320 27807 322 27835
rect 322 27807 354 27835
rect 320 27767 354 27769
rect 320 27735 322 27767
rect 322 27735 354 27767
rect 320 27665 322 27697
rect 322 27665 354 27697
rect 320 27663 354 27665
rect 320 27597 322 27625
rect 322 27597 354 27625
rect 320 27591 354 27597
rect 320 27529 322 27553
rect 322 27529 354 27553
rect 320 27519 354 27529
rect 320 27461 322 27481
rect 322 27461 354 27481
rect 320 27447 354 27461
rect 320 27393 322 27409
rect 322 27393 354 27409
rect 320 27375 354 27393
rect 320 27325 322 27337
rect 322 27325 354 27337
rect 320 27303 354 27325
rect 320 27257 322 27265
rect 322 27257 354 27265
rect 320 27231 354 27257
rect 320 27189 322 27193
rect 322 27189 354 27193
rect 320 27159 354 27189
rect 320 27087 354 27121
rect 320 27019 354 27049
rect 320 27015 322 27019
rect 322 27015 354 27019
rect 320 26951 354 26977
rect 320 26943 322 26951
rect 322 26943 354 26951
rect 320 26883 354 26905
rect 320 26871 322 26883
rect 322 26871 354 26883
rect 320 26815 354 26833
rect 320 26799 322 26815
rect 322 26799 354 26815
rect 320 26747 354 26761
rect 320 26727 322 26747
rect 322 26727 354 26747
rect 320 26679 354 26689
rect 320 26655 322 26679
rect 322 26655 354 26679
rect 320 26611 354 26617
rect 320 26583 322 26611
rect 322 26583 354 26611
rect 320 26543 354 26545
rect 320 26511 322 26543
rect 322 26511 354 26543
rect 320 26441 322 26473
rect 322 26441 354 26473
rect 320 26439 354 26441
rect 320 26373 322 26401
rect 322 26373 354 26401
rect 320 26367 354 26373
rect 320 26305 322 26329
rect 322 26305 354 26329
rect 320 26295 354 26305
rect 320 26237 322 26257
rect 322 26237 354 26257
rect 320 26223 354 26237
rect 320 26169 322 26185
rect 322 26169 354 26185
rect 320 26151 354 26169
rect 320 26101 322 26113
rect 322 26101 354 26113
rect 320 26079 354 26101
rect 320 26033 322 26041
rect 322 26033 354 26041
rect 320 26007 354 26033
rect 320 25965 322 25969
rect 322 25965 354 25969
rect 320 25935 354 25965
rect 320 25863 354 25897
rect 320 25795 354 25825
rect 320 25791 322 25795
rect 322 25791 354 25795
rect 320 25727 354 25753
rect 320 25719 322 25727
rect 322 25719 354 25727
rect 320 25659 354 25681
rect 320 25647 322 25659
rect 322 25647 354 25659
rect 320 25591 354 25609
rect 320 25575 322 25591
rect 322 25575 354 25591
rect 320 25523 354 25537
rect 320 25503 322 25523
rect 322 25503 354 25523
rect 320 25455 354 25465
rect 320 25431 322 25455
rect 322 25431 354 25455
rect 320 25387 354 25393
rect 320 25359 322 25387
rect 322 25359 354 25387
rect 320 25319 354 25321
rect 320 25287 322 25319
rect 322 25287 354 25319
rect 320 25217 322 25249
rect 322 25217 354 25249
rect 320 25215 354 25217
rect 320 25149 322 25177
rect 322 25149 354 25177
rect 320 25143 354 25149
rect 320 25081 322 25105
rect 322 25081 354 25105
rect 320 25071 354 25081
rect 320 25013 322 25033
rect 322 25013 354 25033
rect 320 24999 354 25013
rect 320 24945 322 24961
rect 322 24945 354 24961
rect 320 24927 354 24945
rect 320 24877 322 24889
rect 322 24877 354 24889
rect 320 24855 354 24877
rect 320 24809 322 24817
rect 322 24809 354 24817
rect 320 24783 354 24809
rect 320 24741 322 24745
rect 322 24741 354 24745
rect 320 24711 354 24741
rect 320 24639 354 24673
rect 320 24571 354 24601
rect 320 24567 322 24571
rect 322 24567 354 24571
rect 320 24503 354 24529
rect 320 24495 322 24503
rect 322 24495 354 24503
rect 320 24435 354 24457
rect 320 24423 322 24435
rect 322 24423 354 24435
rect 320 24367 354 24385
rect 320 24351 322 24367
rect 322 24351 354 24367
rect 320 24299 354 24313
rect 320 24279 322 24299
rect 322 24279 354 24299
rect 320 24231 354 24241
rect 320 24207 322 24231
rect 322 24207 354 24231
rect 320 24163 354 24169
rect 320 24135 322 24163
rect 322 24135 354 24163
rect 320 24095 354 24097
rect 320 24063 322 24095
rect 322 24063 354 24095
rect 320 23993 322 24025
rect 322 23993 354 24025
rect 320 23991 354 23993
rect 320 23925 322 23953
rect 322 23925 354 23953
rect 320 23919 354 23925
rect 320 23857 322 23881
rect 322 23857 354 23881
rect 320 23847 354 23857
rect 320 23789 322 23809
rect 322 23789 354 23809
rect 320 23775 354 23789
rect 320 23721 322 23737
rect 322 23721 354 23737
rect 320 23703 354 23721
rect 320 23653 322 23665
rect 322 23653 354 23665
rect 320 23631 354 23653
rect 320 23585 322 23593
rect 322 23585 354 23593
rect 320 23559 354 23585
rect 320 23517 322 23521
rect 322 23517 354 23521
rect 320 23487 354 23517
rect 320 23415 354 23449
rect 320 23347 354 23377
rect 320 23343 322 23347
rect 322 23343 354 23347
rect 320 23279 354 23305
rect 320 23271 322 23279
rect 322 23271 354 23279
rect 320 23211 354 23233
rect 320 23199 322 23211
rect 322 23199 354 23211
rect 320 23143 354 23161
rect 320 23127 322 23143
rect 322 23127 354 23143
rect 320 23075 354 23089
rect 320 23055 322 23075
rect 322 23055 354 23075
rect 320 23007 354 23017
rect 320 22983 322 23007
rect 322 22983 354 23007
rect 320 22939 354 22945
rect 320 22911 322 22939
rect 322 22911 354 22939
rect 320 22871 354 22873
rect 320 22839 322 22871
rect 322 22839 354 22871
rect 320 22769 322 22801
rect 322 22769 354 22801
rect 320 22767 354 22769
rect 320 22701 322 22729
rect 322 22701 354 22729
rect 320 22695 354 22701
rect 320 22633 322 22657
rect 322 22633 354 22657
rect 320 22623 354 22633
rect 320 22565 322 22585
rect 322 22565 354 22585
rect 320 22551 354 22565
rect 320 22497 322 22513
rect 322 22497 354 22513
rect 320 22479 354 22497
rect 320 22429 322 22441
rect 322 22429 354 22441
rect 320 22407 354 22429
rect 320 22361 322 22369
rect 322 22361 354 22369
rect 320 22335 354 22361
rect 320 22293 322 22297
rect 322 22293 354 22297
rect 320 22263 354 22293
rect 320 22191 354 22225
rect 320 22123 354 22153
rect 320 22119 322 22123
rect 322 22119 354 22123
rect 320 22055 354 22081
rect 320 22047 322 22055
rect 322 22047 354 22055
rect 320 21987 354 22009
rect 320 21975 322 21987
rect 322 21975 354 21987
rect 320 21919 354 21937
rect 320 21903 322 21919
rect 322 21903 354 21919
rect 320 21851 354 21865
rect 320 21831 322 21851
rect 322 21831 354 21851
rect 320 21783 354 21793
rect 320 21759 322 21783
rect 322 21759 354 21783
rect 320 21715 354 21721
rect 320 21687 322 21715
rect 322 21687 354 21715
rect 320 21647 354 21649
rect 320 21615 322 21647
rect 322 21615 354 21647
rect 320 21545 322 21577
rect 322 21545 354 21577
rect 320 21543 354 21545
rect 320 21477 322 21505
rect 322 21477 354 21505
rect 320 21471 354 21477
rect 320 21409 322 21433
rect 322 21409 354 21433
rect 320 21399 354 21409
rect 320 21341 322 21361
rect 322 21341 354 21361
rect 320 21327 354 21341
rect 320 21273 322 21289
rect 322 21273 354 21289
rect 320 21255 354 21273
rect 320 21205 322 21217
rect 322 21205 354 21217
rect 320 21183 354 21205
rect 320 21137 322 21145
rect 322 21137 354 21145
rect 320 21111 354 21137
rect 320 21069 322 21073
rect 322 21069 354 21073
rect 320 21039 354 21069
rect 320 20967 354 21001
rect 320 20899 354 20929
rect 320 20895 322 20899
rect 322 20895 354 20899
rect 320 20831 354 20857
rect 320 20823 322 20831
rect 322 20823 354 20831
rect 320 20763 354 20785
rect 320 20751 322 20763
rect 322 20751 354 20763
rect 320 20695 354 20713
rect 320 20679 322 20695
rect 322 20679 354 20695
rect 320 20627 354 20641
rect 320 20607 322 20627
rect 322 20607 354 20627
rect 320 20559 354 20569
rect 320 20535 322 20559
rect 322 20535 354 20559
rect 320 20491 354 20497
rect 320 20463 322 20491
rect 322 20463 354 20491
rect 320 20423 354 20425
rect 320 20391 322 20423
rect 322 20391 354 20423
rect 320 20321 322 20353
rect 322 20321 354 20353
rect 320 20319 354 20321
rect 320 20253 322 20281
rect 322 20253 354 20281
rect 320 20247 354 20253
rect 320 20185 322 20209
rect 322 20185 354 20209
rect 320 20175 354 20185
rect 320 20117 322 20137
rect 322 20117 354 20137
rect 320 20103 354 20117
rect 320 20049 322 20065
rect 322 20049 354 20065
rect 320 20031 354 20049
rect 320 19981 322 19993
rect 322 19981 354 19993
rect 320 19959 354 19981
rect 320 19913 322 19921
rect 322 19913 354 19921
rect 320 19887 354 19913
rect 320 19845 322 19849
rect 322 19845 354 19849
rect 320 19815 354 19845
rect 320 19743 354 19777
rect 320 19675 354 19705
rect 320 19671 322 19675
rect 322 19671 354 19675
rect 320 19607 354 19633
rect 320 19599 322 19607
rect 322 19599 354 19607
rect 320 19539 354 19561
rect 320 19527 322 19539
rect 322 19527 354 19539
rect 320 19471 354 19489
rect 320 19455 322 19471
rect 322 19455 354 19471
rect 320 19403 354 19417
rect 320 19383 322 19403
rect 322 19383 354 19403
rect 320 19335 354 19345
rect 320 19311 322 19335
rect 322 19311 354 19335
rect 320 19267 354 19273
rect 320 19239 322 19267
rect 322 19239 354 19267
rect 320 19199 354 19201
rect 320 19167 322 19199
rect 322 19167 354 19199
rect 320 19097 322 19129
rect 322 19097 354 19129
rect 320 19095 354 19097
rect 320 19029 322 19057
rect 322 19029 354 19057
rect 320 19023 354 19029
rect 320 18961 322 18985
rect 322 18961 354 18985
rect 320 18951 354 18961
rect 320 18893 322 18913
rect 322 18893 354 18913
rect 320 18879 354 18893
rect 320 18825 322 18841
rect 322 18825 354 18841
rect 320 18807 354 18825
rect 320 18757 322 18769
rect 322 18757 354 18769
rect 320 18735 354 18757
rect 320 18689 322 18697
rect 322 18689 354 18697
rect 320 18663 354 18689
rect 320 18621 322 18625
rect 322 18621 354 18625
rect 320 18591 354 18621
rect 320 18519 354 18553
rect 320 18451 354 18481
rect 320 18447 322 18451
rect 322 18447 354 18451
rect 320 18383 354 18409
rect 320 18375 322 18383
rect 322 18375 354 18383
rect 320 18315 354 18337
rect 320 18303 322 18315
rect 322 18303 354 18315
rect 320 18247 354 18265
rect 320 18231 322 18247
rect 322 18231 354 18247
rect 320 18179 354 18193
rect 320 18159 322 18179
rect 322 18159 354 18179
rect 320 18111 354 18121
rect 320 18087 322 18111
rect 322 18087 354 18111
rect 320 18043 354 18049
rect 320 18015 322 18043
rect 322 18015 354 18043
rect 320 17975 354 17977
rect 320 17943 322 17975
rect 322 17943 354 17975
rect 320 17873 322 17905
rect 322 17873 354 17905
rect 320 17871 354 17873
rect 320 17805 322 17833
rect 322 17805 354 17833
rect 320 17799 354 17805
rect 320 17737 322 17761
rect 322 17737 354 17761
rect 320 17727 354 17737
rect 320 17669 322 17689
rect 322 17669 354 17689
rect 320 17655 354 17669
rect 320 17601 322 17617
rect 322 17601 354 17617
rect 320 17583 354 17601
rect 320 17533 322 17545
rect 322 17533 354 17545
rect 320 17511 354 17533
rect 320 17465 322 17473
rect 322 17465 354 17473
rect 320 17439 354 17465
rect 320 17397 322 17401
rect 322 17397 354 17401
rect 320 17367 354 17397
rect 320 17295 354 17329
rect 320 17227 354 17257
rect 320 17223 322 17227
rect 322 17223 354 17227
rect 320 17159 354 17185
rect 320 17151 322 17159
rect 322 17151 354 17159
rect 320 17091 354 17113
rect 320 17079 322 17091
rect 322 17079 354 17091
rect 320 17023 354 17041
rect 320 17007 322 17023
rect 322 17007 354 17023
rect 320 16955 354 16969
rect 320 16935 322 16955
rect 322 16935 354 16955
rect 320 16887 354 16897
rect 320 16863 322 16887
rect 322 16863 354 16887
rect 320 16819 354 16825
rect 320 16791 322 16819
rect 322 16791 354 16819
rect 320 16751 354 16753
rect 320 16719 322 16751
rect 322 16719 354 16751
rect 320 16649 322 16681
rect 322 16649 354 16681
rect 320 16647 354 16649
rect 320 16581 322 16609
rect 322 16581 354 16609
rect 320 16575 354 16581
rect 320 16513 322 16537
rect 322 16513 354 16537
rect 320 16503 354 16513
rect 320 16445 322 16465
rect 322 16445 354 16465
rect 320 16431 354 16445
rect 320 16377 322 16393
rect 322 16377 354 16393
rect 320 16359 354 16377
rect 320 16309 322 16321
rect 322 16309 354 16321
rect 320 16287 354 16309
rect 320 16241 322 16249
rect 322 16241 354 16249
rect 320 16215 354 16241
rect 320 16173 322 16177
rect 322 16173 354 16177
rect 320 16143 354 16173
rect 320 16071 354 16105
rect 320 16003 354 16033
rect 320 15999 322 16003
rect 322 15999 354 16003
rect 320 15935 354 15961
rect 320 15927 322 15935
rect 322 15927 354 15935
rect 320 15867 354 15889
rect 320 15855 322 15867
rect 322 15855 354 15867
rect 320 15799 354 15817
rect 320 15783 322 15799
rect 322 15783 354 15799
rect 320 15731 354 15745
rect 320 15711 322 15731
rect 322 15711 354 15731
rect 320 15663 354 15673
rect 320 15639 322 15663
rect 322 15639 354 15663
rect 320 15595 354 15601
rect 320 15567 322 15595
rect 322 15567 354 15595
rect 320 15527 354 15529
rect 320 15495 322 15527
rect 322 15495 354 15527
rect 320 15425 322 15457
rect 322 15425 354 15457
rect 320 15423 354 15425
rect 320 15357 322 15385
rect 322 15357 354 15385
rect 320 15351 354 15357
rect 320 15289 322 15313
rect 322 15289 354 15313
rect 320 15279 354 15289
rect 320 15221 322 15241
rect 322 15221 354 15241
rect 320 15207 354 15221
rect 320 15153 322 15169
rect 322 15153 354 15169
rect 320 15135 354 15153
rect 320 15085 322 15097
rect 322 15085 354 15097
rect 320 15063 354 15085
rect 320 15017 322 15025
rect 322 15017 354 15025
rect 320 14991 354 15017
rect 320 14949 322 14953
rect 322 14949 354 14953
rect 320 14919 354 14949
rect 320 14847 354 14881
rect 320 14779 354 14809
rect 320 14775 322 14779
rect 322 14775 354 14779
rect 320 14711 354 14737
rect 320 14703 322 14711
rect 322 14703 354 14711
rect 320 14643 354 14665
rect 320 14631 322 14643
rect 322 14631 354 14643
rect 320 14575 354 14593
rect 320 14559 322 14575
rect 322 14559 354 14575
rect 320 14507 354 14521
rect 320 14487 322 14507
rect 322 14487 354 14507
rect 320 14439 354 14449
rect 320 14415 322 14439
rect 322 14415 354 14439
rect 320 14371 354 14377
rect 320 14343 322 14371
rect 322 14343 354 14371
rect 320 14303 354 14305
rect 320 14271 322 14303
rect 322 14271 354 14303
rect 320 14201 322 14233
rect 322 14201 354 14233
rect 320 14199 354 14201
rect 320 14133 322 14161
rect 322 14133 354 14161
rect 320 14127 354 14133
rect 320 14065 322 14089
rect 322 14065 354 14089
rect 320 14055 354 14065
rect 320 13997 322 14017
rect 322 13997 354 14017
rect 320 13983 354 13997
rect 320 13929 322 13945
rect 322 13929 354 13945
rect 320 13911 354 13929
rect 320 13861 322 13873
rect 322 13861 354 13873
rect 320 13839 354 13861
rect 320 13793 322 13801
rect 322 13793 354 13801
rect 320 13767 354 13793
rect 320 13725 322 13729
rect 322 13725 354 13729
rect 320 13695 354 13725
rect 320 13623 354 13657
rect 320 13555 354 13585
rect 320 13551 322 13555
rect 322 13551 354 13555
rect 320 13487 354 13513
rect 320 13479 322 13487
rect 322 13479 354 13487
rect 320 13419 354 13441
rect 320 13407 322 13419
rect 322 13407 354 13419
rect 320 13351 354 13369
rect 320 13335 322 13351
rect 322 13335 354 13351
rect 320 13283 354 13297
rect 320 13263 322 13283
rect 322 13263 354 13283
rect 320 13215 354 13225
rect 320 13191 322 13215
rect 322 13191 354 13215
rect 320 13147 354 13153
rect 320 13119 322 13147
rect 322 13119 354 13147
rect 320 13079 354 13081
rect 320 13047 322 13079
rect 322 13047 354 13079
rect 320 12977 322 13009
rect 322 12977 354 13009
rect 320 12975 354 12977
rect 320 12909 322 12937
rect 322 12909 354 12937
rect 320 12903 354 12909
rect 320 12841 322 12865
rect 322 12841 354 12865
rect 320 12831 354 12841
rect 320 12773 322 12793
rect 322 12773 354 12793
rect 320 12759 354 12773
rect 320 12705 322 12721
rect 322 12705 354 12721
rect 320 12687 354 12705
rect 320 12637 322 12649
rect 322 12637 354 12649
rect 320 12615 354 12637
rect 320 12569 322 12577
rect 322 12569 354 12577
rect 320 12543 354 12569
rect 320 12501 322 12505
rect 322 12501 354 12505
rect 320 12471 354 12501
rect 320 12399 354 12433
rect 320 12331 354 12361
rect 320 12327 322 12331
rect 322 12327 354 12331
rect 320 12263 354 12289
rect 320 12255 322 12263
rect 322 12255 354 12263
rect 320 12195 354 12217
rect 320 12183 322 12195
rect 322 12183 354 12195
rect 320 12127 354 12145
rect 320 12111 322 12127
rect 322 12111 354 12127
rect 320 12059 354 12073
rect 320 12039 322 12059
rect 322 12039 354 12059
rect 320 11991 354 12001
rect 320 11967 322 11991
rect 322 11967 354 11991
rect 320 11923 354 11929
rect 320 11895 322 11923
rect 322 11895 354 11923
rect 320 11855 354 11857
rect 320 11823 322 11855
rect 322 11823 354 11855
rect 320 11753 322 11785
rect 322 11753 354 11785
rect 320 11751 354 11753
rect 320 11685 322 11713
rect 322 11685 354 11713
rect 320 11679 354 11685
rect 320 11617 322 11641
rect 322 11617 354 11641
rect 320 11607 354 11617
rect 320 11549 322 11569
rect 322 11549 354 11569
rect 320 11535 354 11549
rect 320 11481 322 11497
rect 322 11481 354 11497
rect 320 11463 354 11481
rect 320 11413 322 11425
rect 322 11413 354 11425
rect 320 11391 354 11413
rect 320 11345 322 11353
rect 322 11345 354 11353
rect 320 11319 354 11345
rect 320 11277 322 11281
rect 322 11277 354 11281
rect 320 11247 354 11277
rect 320 11175 354 11209
rect 320 11107 354 11137
rect 320 11103 322 11107
rect 322 11103 354 11107
rect 320 11039 354 11065
rect 320 11031 322 11039
rect 322 11031 354 11039
rect 320 10971 354 10993
rect 320 10959 322 10971
rect 322 10959 354 10971
rect 320 10903 354 10921
rect 320 10887 322 10903
rect 322 10887 354 10903
rect 320 10835 354 10849
rect 320 10815 322 10835
rect 322 10815 354 10835
rect 320 10767 354 10777
rect 320 10743 322 10767
rect 322 10743 354 10767
rect 320 10699 354 10705
rect 320 10671 322 10699
rect 322 10671 354 10699
rect 320 10631 354 10633
rect 320 10599 322 10631
rect 322 10599 354 10631
rect 320 10529 322 10561
rect 322 10529 354 10561
rect 320 10527 354 10529
rect 320 10461 322 10489
rect 322 10461 354 10489
rect 320 10455 354 10461
rect 320 10393 322 10417
rect 322 10393 354 10417
rect 320 10383 354 10393
rect 320 10325 322 10345
rect 322 10325 354 10345
rect 320 10311 354 10325
rect 320 10257 322 10273
rect 322 10257 354 10273
rect 320 10239 354 10257
rect 320 10189 322 10201
rect 322 10189 354 10201
rect 320 10167 354 10189
rect 320 10121 322 10129
rect 322 10121 354 10129
rect 320 10095 354 10121
rect 320 10053 322 10057
rect 322 10053 354 10057
rect 320 10023 354 10053
rect 320 9951 354 9985
rect 320 9883 354 9913
rect 320 9879 322 9883
rect 322 9879 354 9883
rect 320 9815 354 9841
rect 320 9807 322 9815
rect 322 9807 354 9815
rect 320 9747 354 9769
rect 320 9735 322 9747
rect 322 9735 354 9747
rect 1009 35969 1043 36003
rect 1081 35969 1115 36003
rect 1153 35969 1187 36003
rect 1225 35969 1259 36003
rect 1297 35969 1331 36003
rect 1369 35969 1403 36003
rect 1441 35969 1475 36003
rect 1513 35969 1547 36003
rect 1585 35969 1619 36003
rect 1657 35969 1691 36003
rect 1729 35969 1763 36003
rect 1801 35969 1835 36003
rect 1873 35969 1907 36003
rect 1945 35969 1979 36003
rect 2017 35969 2051 36003
rect 2089 35969 2123 36003
rect 2161 35969 2195 36003
rect 2233 35969 2267 36003
rect 2305 35969 2339 36003
rect 2377 35969 2411 36003
rect 2449 35969 2483 36003
rect 2521 35969 2555 36003
rect 2593 35969 2627 36003
rect 2665 35969 2699 36003
rect 2737 35969 2771 36003
rect 2809 35969 2843 36003
rect 2881 35969 2915 36003
rect 2953 35969 2987 36003
rect 3025 35969 3059 36003
rect 3097 35969 3131 36003
rect 3169 35969 3203 36003
rect 3241 35969 3275 36003
rect 3313 35969 3347 36003
rect 3385 35969 3419 36003
rect 3457 35969 3491 36003
rect 3529 35969 3563 36003
rect 3601 35969 3635 36003
rect 3673 35969 3707 36003
rect 3745 35969 3779 36003
rect 3817 35969 3851 36003
rect 3889 35969 3923 36003
rect 3961 35969 3995 36003
rect 4033 35969 4067 36003
rect 4105 35969 4139 36003
rect 4177 35969 4211 36003
rect 4249 35969 4283 36003
rect 4321 35969 4355 36003
rect 4393 35969 4427 36003
rect 4465 35969 4499 36003
rect 4537 35969 4571 36003
rect 4609 35969 4643 36003
rect 4681 35969 4715 36003
rect 4753 35969 4787 36003
rect 4825 35969 4859 36003
rect 4897 35969 4931 36003
rect 4969 35969 5003 36003
rect 5041 35969 5075 36003
rect 5113 35969 5147 36003
rect 5185 35969 5219 36003
rect 5257 35969 5291 36003
rect 5329 35969 5363 36003
rect 5401 35969 5435 36003
rect 5473 35969 5507 36003
rect 5545 35969 5579 36003
rect 5617 35969 5651 36003
rect 5689 35969 5723 36003
rect 5761 35969 5795 36003
rect 5833 35969 5867 36003
rect 5905 35969 5939 36003
rect 5977 35969 6011 36003
rect 6049 35969 6083 36003
rect 6121 35969 6155 36003
rect 6193 35969 6227 36003
rect 6265 35969 6299 36003
rect 6337 35969 6371 36003
rect 6409 35969 6443 36003
rect 6481 35969 6515 36003
rect 6553 35969 6587 36003
rect 6625 35969 6659 36003
rect 6697 35969 6731 36003
rect 6769 35969 6803 36003
rect 6841 35969 6875 36003
rect 6913 35969 6947 36003
rect 6985 35969 7019 36003
rect 7057 35969 7091 36003
rect 7129 35969 7163 36003
rect 7201 35969 7235 36003
rect 7273 35969 7307 36003
rect 7345 35969 7379 36003
rect 7417 35969 7451 36003
rect 7489 35969 7523 36003
rect 7561 35969 7595 36003
rect 7633 35969 7667 36003
rect 7705 35969 7739 36003
rect 7777 35969 7811 36003
rect 7849 35969 7883 36003
rect 7921 35969 7955 36003
rect 7993 35969 8027 36003
rect 8065 35969 8099 36003
rect 8137 35969 8171 36003
rect 8209 35969 8243 36003
rect 8281 35969 8315 36003
rect 8353 35969 8387 36003
rect 8425 35969 8459 36003
rect 8497 35969 8531 36003
rect 8569 35969 8603 36003
rect 8641 35969 8675 36003
rect 8713 35969 8747 36003
rect 8785 35969 8819 36003
rect 8857 35969 8891 36003
rect 8929 35969 8963 36003
rect 9001 35969 9035 36003
rect 9073 35969 9107 36003
rect 9145 35969 9179 36003
rect 9217 35969 9251 36003
rect 9289 35969 9323 36003
rect 9361 35969 9395 36003
rect 9433 35969 9467 36003
rect 9505 35969 9539 36003
rect 9577 35969 9611 36003
rect 9649 35969 9683 36003
rect 9721 35969 9755 36003
rect 9793 35969 9827 36003
rect 9865 35969 9899 36003
rect 9937 35969 9971 36003
rect 10009 35969 10043 36003
rect 10081 35969 10115 36003
rect 10153 35969 10187 36003
rect 10225 35969 10259 36003
rect 10297 35969 10331 36003
rect 10369 35969 10403 36003
rect 10441 35969 10475 36003
rect 10513 35969 10547 36003
rect 10585 35969 10619 36003
rect 10657 35969 10691 36003
rect 10729 35969 10763 36003
rect 10801 35969 10835 36003
rect 10873 35969 10907 36003
rect 10945 35969 10979 36003
rect 11017 35969 11051 36003
rect 11089 35969 11123 36003
rect 11161 35969 11195 36003
rect 11233 35969 11267 36003
rect 11305 35969 11339 36003
rect 11377 35969 11411 36003
rect 11449 35969 11483 36003
rect 11521 35969 11555 36003
rect 11593 35969 11627 36003
rect 11665 35969 11699 36003
rect 11737 35969 11771 36003
rect 11809 35969 11843 36003
rect 11881 35969 11915 36003
rect 11953 35969 11987 36003
rect 12025 35969 12059 36003
rect 12097 35969 12131 36003
rect 12169 35969 12203 36003
rect 12241 35969 12275 36003
rect 12313 35969 12347 36003
rect 12385 35969 12419 36003
rect 12457 35969 12491 36003
rect 12529 35969 12563 36003
rect 12601 35969 12635 36003
rect 12673 35969 12707 36003
rect 12745 35969 12779 36003
rect 12817 35969 12851 36003
rect 12889 35969 12923 36003
rect 12961 35969 12995 36003
rect 13033 35969 13067 36003
rect 13105 35969 13139 36003
rect 13177 35969 13211 36003
rect 13249 35969 13283 36003
rect 13321 35969 13355 36003
rect 13393 35969 13427 36003
rect 13465 35969 13499 36003
rect 13537 35969 13571 36003
rect 13609 35969 13643 36003
rect 13681 35969 13715 36003
rect 13753 35969 13787 36003
rect 13825 35969 13859 36003
rect 13897 35969 13931 36003
rect 13969 35969 14003 36003
rect 814 35877 848 35911
rect 814 35805 848 35839
rect 14120 35798 14154 35832
rect 814 35733 848 35767
rect 14120 35726 14154 35760
rect 814 35661 848 35695
rect 14120 35654 14154 35688
rect 814 35589 848 35623
rect 14120 35582 14154 35616
rect 814 35517 848 35551
rect 14120 35510 14154 35544
rect 814 35445 848 35479
rect 14120 35438 14154 35472
rect 814 35373 848 35407
rect 14120 35366 14154 35400
rect 814 35301 848 35335
rect 14120 35294 14154 35328
rect 814 35229 848 35263
rect 14120 35222 14154 35256
rect 814 35157 848 35191
rect 14120 35150 14154 35184
rect 814 35085 848 35119
rect 14120 35078 14154 35112
rect 814 35013 848 35047
rect 14120 35006 14154 35040
rect 814 34941 848 34975
rect 14120 34934 14154 34968
rect 814 34869 848 34903
rect 14120 34862 14154 34896
rect 814 34797 848 34831
rect 814 34725 848 34759
rect 814 34653 848 34687
rect 14120 34790 14154 34824
rect 14120 34718 14154 34752
rect 814 34581 848 34615
rect 814 34509 848 34543
rect 814 34437 848 34471
rect 814 34365 848 34399
rect 814 34293 848 34327
rect 814 34221 848 34255
rect 814 34149 848 34183
rect 814 34077 848 34111
rect 814 34005 848 34039
rect 814 33933 848 33967
rect 814 33861 848 33895
rect 814 33789 848 33823
rect 814 33717 848 33751
rect 814 33645 848 33679
rect 814 33573 848 33607
rect 814 33501 848 33535
rect 814 33429 848 33463
rect 814 33357 848 33391
rect 814 33285 848 33319
rect 814 33213 848 33247
rect 814 33141 848 33175
rect 814 33069 848 33103
rect 814 32997 848 33031
rect 814 32925 848 32959
rect 814 32853 848 32887
rect 814 32781 848 32815
rect 814 32709 848 32743
rect 814 32637 848 32671
rect 814 32565 848 32599
rect 814 32493 848 32527
rect 814 32421 848 32455
rect 814 32349 848 32383
rect 814 32277 848 32311
rect 814 32205 848 32239
rect 814 32133 848 32167
rect 814 32061 848 32095
rect 814 31989 848 32023
rect 814 31917 848 31951
rect 814 31845 848 31879
rect 814 31773 848 31807
rect 814 31701 848 31735
rect 814 31629 848 31663
rect 814 31557 848 31591
rect 814 31485 848 31519
rect 814 31413 848 31447
rect 814 31341 848 31375
rect 814 31269 848 31303
rect 814 31197 848 31231
rect 814 31125 848 31159
rect 814 31053 848 31087
rect 814 30981 848 31015
rect 814 30909 848 30943
rect 814 30837 848 30871
rect 814 30765 848 30799
rect 814 30693 848 30727
rect 814 30621 848 30655
rect 814 30549 848 30583
rect 814 30477 848 30511
rect 814 30405 848 30439
rect 814 30333 848 30367
rect 814 30261 848 30295
rect 814 30189 848 30223
rect 814 30117 848 30151
rect 814 30045 848 30079
rect 814 29973 848 30007
rect 814 29901 848 29935
rect 814 29829 848 29863
rect 814 29757 848 29791
rect 814 29685 848 29719
rect 814 29613 848 29647
rect 814 29541 848 29575
rect 814 29469 848 29503
rect 814 29397 848 29431
rect 814 29325 848 29359
rect 814 29253 848 29287
rect 814 29181 848 29215
rect 814 29109 848 29143
rect 814 29037 848 29071
rect 814 28965 848 28999
rect 814 28893 848 28927
rect 814 28821 848 28855
rect 814 28749 848 28783
rect 814 28677 848 28711
rect 814 28605 848 28639
rect 814 28533 848 28567
rect 814 28461 848 28495
rect 814 28389 848 28423
rect 814 28317 848 28351
rect 814 28245 848 28279
rect 814 28173 848 28207
rect 814 28101 848 28135
rect 814 28029 848 28063
rect 814 27957 848 27991
rect 814 27885 848 27919
rect 814 27813 848 27847
rect 814 27741 848 27775
rect 814 27669 848 27703
rect 814 27597 848 27631
rect 814 27525 848 27559
rect 814 27453 848 27487
rect 814 27381 848 27415
rect 814 27309 848 27343
rect 814 27237 848 27271
rect 814 27165 848 27199
rect 814 27093 848 27127
rect 814 27021 848 27055
rect 814 26949 848 26983
rect 814 26877 848 26911
rect 814 26805 848 26839
rect 814 26733 848 26767
rect 814 26661 848 26695
rect 814 26589 848 26623
rect 814 26517 848 26551
rect 814 26445 848 26479
rect 814 26373 848 26407
rect 814 26301 848 26335
rect 814 26229 848 26263
rect 814 26157 848 26191
rect 814 26085 848 26119
rect 814 26013 848 26047
rect 814 25941 848 25975
rect 814 25869 848 25903
rect 814 25797 848 25831
rect 814 25725 848 25759
rect 814 25653 848 25687
rect 814 25581 848 25615
rect 814 25509 848 25543
rect 814 25437 848 25471
rect 814 25365 848 25399
rect 814 25293 848 25327
rect 814 25221 848 25255
rect 814 25149 848 25183
rect 814 25077 848 25111
rect 814 25005 848 25039
rect 814 24933 848 24967
rect 814 24861 848 24895
rect 814 24789 848 24823
rect 814 24717 848 24751
rect 814 24645 848 24679
rect 814 24573 848 24607
rect 814 24501 848 24535
rect 814 24429 848 24463
rect 814 24357 848 24391
rect 814 24285 848 24319
rect 814 24213 848 24247
rect 814 24141 848 24175
rect 814 24069 848 24103
rect 814 23997 848 24031
rect 814 23925 848 23959
rect 814 23853 848 23887
rect 814 23781 848 23815
rect 814 23709 848 23743
rect 814 23637 848 23671
rect 814 23565 848 23599
rect 814 23493 848 23527
rect 814 23421 848 23455
rect 814 23349 848 23383
rect 814 23277 848 23311
rect 814 23205 848 23239
rect 814 23133 848 23167
rect 814 23061 848 23095
rect 814 22989 848 23023
rect 814 22917 848 22951
rect 814 22845 848 22879
rect 814 22773 848 22807
rect 814 22701 848 22735
rect 814 22629 848 22663
rect 814 22557 848 22591
rect 814 22485 848 22519
rect 814 22413 848 22447
rect 814 22341 848 22375
rect 814 22269 848 22303
rect 814 22197 848 22231
rect 814 22125 848 22159
rect 814 22053 848 22087
rect 814 21981 848 22015
rect 814 21909 848 21943
rect 814 21837 848 21871
rect 814 21765 848 21799
rect 814 21693 848 21727
rect 814 21621 848 21655
rect 814 21549 848 21583
rect 814 21477 848 21511
rect 814 21405 848 21439
rect 814 21333 848 21367
rect 814 21261 848 21295
rect 814 21189 848 21223
rect 814 21117 848 21151
rect 814 21045 848 21079
rect 814 20973 848 21007
rect 814 20901 848 20935
rect 814 20829 848 20863
rect 814 20757 848 20791
rect 814 20685 848 20719
rect 814 20613 848 20647
rect 814 20541 848 20575
rect 814 20469 848 20503
rect 814 20397 848 20431
rect 814 20325 848 20359
rect 814 20253 848 20287
rect 814 20181 848 20215
rect 814 20109 848 20143
rect 814 20037 848 20071
rect 814 19965 848 19999
rect 814 19893 848 19927
rect 814 19821 848 19855
rect 814 19749 848 19783
rect 814 19677 848 19711
rect 814 19605 848 19639
rect 814 19533 848 19567
rect 814 19461 848 19495
rect 814 19389 848 19423
rect 814 19317 848 19351
rect 814 19245 848 19279
rect 814 19173 848 19207
rect 814 19101 848 19135
rect 814 19029 848 19063
rect 814 18957 848 18991
rect 814 18885 848 18919
rect 814 18813 848 18847
rect 814 18741 848 18775
rect 814 18669 848 18703
rect 814 18597 848 18631
rect 814 18525 848 18559
rect 814 18453 848 18487
rect 814 18381 848 18415
rect 814 18309 848 18343
rect 814 18237 848 18271
rect 814 18165 848 18199
rect 814 18093 848 18127
rect 814 18021 848 18055
rect 814 17949 848 17983
rect 814 17877 848 17911
rect 814 17805 848 17839
rect 814 17733 848 17767
rect 814 17661 848 17695
rect 814 17589 848 17623
rect 814 17517 848 17551
rect 814 17445 848 17479
rect 814 17373 848 17407
rect 814 17301 848 17335
rect 814 17229 848 17263
rect 814 17157 848 17191
rect 814 17085 848 17119
rect 814 17013 848 17047
rect 814 16941 848 16975
rect 814 16869 848 16903
rect 814 16797 848 16831
rect 814 16725 848 16759
rect 814 16653 848 16687
rect 814 16581 848 16615
rect 814 16509 848 16543
rect 814 16437 848 16471
rect 814 16365 848 16399
rect 814 16293 848 16327
rect 814 16221 848 16255
rect 814 16149 848 16183
rect 814 16077 848 16111
rect 814 16005 848 16039
rect 814 15933 848 15967
rect 814 15861 848 15895
rect 814 15789 848 15823
rect 814 15717 848 15751
rect 814 15645 848 15679
rect 814 15573 848 15607
rect 814 15501 848 15535
rect 814 15429 848 15463
rect 814 15357 848 15391
rect 814 15285 848 15319
rect 814 15213 848 15247
rect 814 15141 848 15175
rect 814 15069 848 15103
rect 814 14997 848 15031
rect 814 14925 848 14959
rect 814 14853 848 14887
rect 814 14781 848 14815
rect 814 14709 848 14743
rect 814 14637 848 14671
rect 814 14565 848 14599
rect 814 14493 848 14527
rect 814 14421 848 14455
rect 814 14349 848 14383
rect 814 14277 848 14311
rect 814 14205 848 14239
rect 814 14133 848 14167
rect 814 14061 848 14095
rect 814 13989 848 14023
rect 814 13917 848 13951
rect 814 13845 848 13879
rect 814 13773 848 13807
rect 814 13701 848 13735
rect 814 13629 848 13663
rect 814 13557 848 13591
rect 814 13485 848 13519
rect 814 13413 848 13447
rect 814 13341 848 13375
rect 814 13269 848 13303
rect 814 13197 848 13231
rect 814 13125 848 13159
rect 814 13053 848 13087
rect 814 12981 848 13015
rect 814 12909 848 12943
rect 814 12837 848 12871
rect 814 12765 848 12799
rect 814 12693 848 12727
rect 814 12621 848 12655
rect 814 12549 848 12583
rect 814 12477 848 12511
rect 814 12405 848 12439
rect 814 12333 848 12367
rect 814 12261 848 12295
rect 814 12189 848 12223
rect 814 12117 848 12151
rect 814 12045 848 12079
rect 814 11973 848 12007
rect 814 11901 848 11935
rect 814 11829 848 11863
rect 814 11757 848 11791
rect 814 11685 848 11719
rect 814 11613 848 11647
rect 814 11541 848 11575
rect 814 11469 848 11503
rect 814 11397 848 11431
rect 814 11325 848 11359
rect 814 11253 848 11287
rect 814 11181 848 11215
rect 814 11109 848 11143
rect 814 11037 848 11071
rect 814 10965 848 10999
rect 814 10893 848 10927
rect 814 10821 848 10855
rect 814 10749 848 10783
rect 814 10677 848 10711
rect 814 10605 848 10639
rect 814 10533 848 10567
rect 814 10461 848 10495
rect 814 10389 848 10423
rect 814 10317 848 10351
rect 814 10245 848 10279
rect 1365 34602 1399 34636
rect 1437 34602 1467 34636
rect 1467 34602 1471 34636
rect 1509 34602 1535 34636
rect 1535 34602 1543 34636
rect 1581 34602 1603 34636
rect 1603 34602 1615 34636
rect 1653 34602 1671 34636
rect 1671 34602 1687 34636
rect 1725 34602 1739 34636
rect 1739 34602 1759 34636
rect 1797 34602 1807 34636
rect 1807 34602 1831 34636
rect 1869 34602 1875 34636
rect 1875 34602 1903 34636
rect 1941 34602 1943 34636
rect 1943 34602 1975 34636
rect 2013 34602 2045 34636
rect 2045 34602 2047 34636
rect 2085 34602 2113 34636
rect 2113 34602 2119 34636
rect 2157 34602 2181 34636
rect 2181 34602 2191 34636
rect 2229 34602 2249 34636
rect 2249 34602 2263 34636
rect 2301 34602 2317 34636
rect 2317 34602 2335 34636
rect 2373 34602 2385 34636
rect 2385 34602 2407 34636
rect 2445 34602 2453 34636
rect 2453 34602 2479 34636
rect 2517 34602 2521 34636
rect 2521 34602 2551 34636
rect 2589 34602 2623 34636
rect 2661 34602 2691 34636
rect 2691 34602 2695 34636
rect 2733 34602 2759 34636
rect 2759 34602 2767 34636
rect 2805 34602 2827 34636
rect 2827 34602 2839 34636
rect 2877 34602 2895 34636
rect 2895 34602 2911 34636
rect 2949 34602 2963 34636
rect 2963 34602 2983 34636
rect 3021 34602 3031 34636
rect 3031 34602 3055 34636
rect 3093 34602 3099 34636
rect 3099 34602 3127 34636
rect 3165 34602 3167 34636
rect 3167 34602 3199 34636
rect 3237 34602 3269 34636
rect 3269 34602 3271 34636
rect 3309 34602 3337 34636
rect 3337 34602 3343 34636
rect 3381 34602 3405 34636
rect 3405 34602 3415 34636
rect 3453 34602 3473 34636
rect 3473 34602 3487 34636
rect 3525 34602 3541 34636
rect 3541 34602 3559 34636
rect 3597 34602 3609 34636
rect 3609 34602 3631 34636
rect 3669 34602 3677 34636
rect 3677 34602 3703 34636
rect 3741 34602 3745 34636
rect 3745 34602 3775 34636
rect 3813 34602 3847 34636
rect 3885 34602 3915 34636
rect 3915 34602 3919 34636
rect 3957 34602 3983 34636
rect 3983 34602 3991 34636
rect 4029 34602 4051 34636
rect 4051 34602 4063 34636
rect 4101 34602 4119 34636
rect 4119 34602 4135 34636
rect 4173 34602 4187 34636
rect 4187 34602 4207 34636
rect 4245 34602 4255 34636
rect 4255 34602 4279 34636
rect 4317 34602 4323 34636
rect 4323 34602 4351 34636
rect 4389 34602 4391 34636
rect 4391 34602 4423 34636
rect 4461 34602 4493 34636
rect 4493 34602 4495 34636
rect 4533 34602 4561 34636
rect 4561 34602 4567 34636
rect 4605 34602 4629 34636
rect 4629 34602 4639 34636
rect 4677 34602 4697 34636
rect 4697 34602 4711 34636
rect 4749 34602 4765 34636
rect 4765 34602 4783 34636
rect 4821 34602 4833 34636
rect 4833 34602 4855 34636
rect 4893 34602 4901 34636
rect 4901 34602 4927 34636
rect 4965 34602 4969 34636
rect 4969 34602 4999 34636
rect 5037 34602 5071 34636
rect 5109 34602 5139 34636
rect 5139 34602 5143 34636
rect 5181 34602 5207 34636
rect 5207 34602 5215 34636
rect 5253 34602 5275 34636
rect 5275 34602 5287 34636
rect 5325 34602 5343 34636
rect 5343 34602 5359 34636
rect 5397 34602 5411 34636
rect 5411 34602 5431 34636
rect 5469 34602 5479 34636
rect 5479 34602 5503 34636
rect 5541 34602 5547 34636
rect 5547 34602 5575 34636
rect 5613 34602 5615 34636
rect 5615 34602 5647 34636
rect 5685 34602 5717 34636
rect 5717 34602 5719 34636
rect 5757 34602 5785 34636
rect 5785 34602 5791 34636
rect 5829 34602 5853 34636
rect 5853 34602 5863 34636
rect 5901 34602 5921 34636
rect 5921 34602 5935 34636
rect 5973 34602 5989 34636
rect 5989 34602 6007 34636
rect 6045 34602 6057 34636
rect 6057 34602 6079 34636
rect 6117 34602 6125 34636
rect 6125 34602 6151 34636
rect 6189 34602 6193 34636
rect 6193 34602 6223 34636
rect 6261 34602 6295 34636
rect 6333 34602 6363 34636
rect 6363 34602 6367 34636
rect 6405 34602 6431 34636
rect 6431 34602 6439 34636
rect 6477 34602 6499 34636
rect 6499 34602 6511 34636
rect 6549 34602 6567 34636
rect 6567 34602 6583 34636
rect 6621 34602 6635 34636
rect 6635 34602 6655 34636
rect 6693 34602 6703 34636
rect 6703 34602 6727 34636
rect 6765 34602 6771 34636
rect 6771 34602 6799 34636
rect 6837 34602 6839 34636
rect 6839 34602 6871 34636
rect 6909 34602 6941 34636
rect 6941 34602 6943 34636
rect 6981 34602 7009 34636
rect 7009 34602 7015 34636
rect 7053 34602 7077 34636
rect 7077 34602 7087 34636
rect 7125 34602 7145 34636
rect 7145 34602 7159 34636
rect 7197 34602 7213 34636
rect 7213 34602 7231 34636
rect 7269 34602 7281 34636
rect 7281 34602 7303 34636
rect 7341 34602 7349 34636
rect 7349 34602 7375 34636
rect 7413 34602 7417 34636
rect 7417 34602 7447 34636
rect 7485 34602 7519 34636
rect 7557 34602 7587 34636
rect 7587 34602 7591 34636
rect 7629 34602 7655 34636
rect 7655 34602 7663 34636
rect 7701 34602 7723 34636
rect 7723 34602 7735 34636
rect 7773 34602 7791 34636
rect 7791 34602 7807 34636
rect 7845 34602 7859 34636
rect 7859 34602 7879 34636
rect 7917 34602 7927 34636
rect 7927 34602 7951 34636
rect 7989 34602 7995 34636
rect 7995 34602 8023 34636
rect 8061 34602 8063 34636
rect 8063 34602 8095 34636
rect 8133 34602 8165 34636
rect 8165 34602 8167 34636
rect 8205 34602 8233 34636
rect 8233 34602 8239 34636
rect 8277 34602 8301 34636
rect 8301 34602 8311 34636
rect 8349 34602 8369 34636
rect 8369 34602 8383 34636
rect 8421 34602 8437 34636
rect 8437 34602 8455 34636
rect 8493 34602 8505 34636
rect 8505 34602 8527 34636
rect 8565 34602 8573 34636
rect 8573 34602 8599 34636
rect 8637 34602 8641 34636
rect 8641 34602 8671 34636
rect 8709 34602 8743 34636
rect 8781 34602 8811 34636
rect 8811 34602 8815 34636
rect 8853 34602 8879 34636
rect 8879 34602 8887 34636
rect 8925 34602 8947 34636
rect 8947 34602 8959 34636
rect 8997 34602 9015 34636
rect 9015 34602 9031 34636
rect 9069 34602 9083 34636
rect 9083 34602 9103 34636
rect 9141 34602 9151 34636
rect 9151 34602 9175 34636
rect 9213 34602 9219 34636
rect 9219 34602 9247 34636
rect 9285 34602 9287 34636
rect 9287 34602 9319 34636
rect 9357 34602 9389 34636
rect 9389 34602 9391 34636
rect 9429 34602 9457 34636
rect 9457 34602 9463 34636
rect 9501 34602 9525 34636
rect 9525 34602 9535 34636
rect 9573 34602 9593 34636
rect 9593 34602 9607 34636
rect 9645 34602 9661 34636
rect 9661 34602 9679 34636
rect 9717 34602 9729 34636
rect 9729 34602 9751 34636
rect 9789 34602 9797 34636
rect 9797 34602 9823 34636
rect 9861 34602 9865 34636
rect 9865 34602 9895 34636
rect 9933 34602 9967 34636
rect 10005 34602 10035 34636
rect 10035 34602 10039 34636
rect 10077 34602 10103 34636
rect 10103 34602 10111 34636
rect 10149 34602 10171 34636
rect 10171 34602 10183 34636
rect 10221 34602 10239 34636
rect 10239 34602 10255 34636
rect 10293 34602 10307 34636
rect 10307 34602 10327 34636
rect 10365 34602 10375 34636
rect 10375 34602 10399 34636
rect 10437 34602 10443 34636
rect 10443 34602 10471 34636
rect 10509 34602 10511 34636
rect 10511 34602 10543 34636
rect 10581 34602 10613 34636
rect 10613 34602 10615 34636
rect 10653 34602 10681 34636
rect 10681 34602 10687 34636
rect 10725 34602 10749 34636
rect 10749 34602 10759 34636
rect 10797 34602 10817 34636
rect 10817 34602 10831 34636
rect 10869 34602 10885 34636
rect 10885 34602 10903 34636
rect 10941 34602 10953 34636
rect 10953 34602 10975 34636
rect 11013 34602 11021 34636
rect 11021 34602 11047 34636
rect 11085 34602 11089 34636
rect 11089 34602 11119 34636
rect 11157 34602 11191 34636
rect 11229 34602 11259 34636
rect 11259 34602 11263 34636
rect 11301 34602 11327 34636
rect 11327 34602 11335 34636
rect 11373 34602 11395 34636
rect 11395 34602 11407 34636
rect 11445 34602 11463 34636
rect 11463 34602 11479 34636
rect 11517 34602 11531 34636
rect 11531 34602 11551 34636
rect 11589 34602 11599 34636
rect 11599 34602 11623 34636
rect 11661 34602 11667 34636
rect 11667 34602 11695 34636
rect 11733 34602 11735 34636
rect 11735 34602 11767 34636
rect 11805 34602 11837 34636
rect 11837 34602 11839 34636
rect 11877 34602 11905 34636
rect 11905 34602 11911 34636
rect 11949 34602 11973 34636
rect 11973 34602 11983 34636
rect 12021 34602 12041 34636
rect 12041 34602 12055 34636
rect 12093 34602 12109 34636
rect 12109 34602 12127 34636
rect 12165 34602 12177 34636
rect 12177 34602 12199 34636
rect 12237 34602 12245 34636
rect 12245 34602 12271 34636
rect 12309 34602 12313 34636
rect 12313 34602 12343 34636
rect 12381 34602 12415 34636
rect 12453 34602 12483 34636
rect 12483 34602 12487 34636
rect 12525 34602 12551 34636
rect 12551 34602 12559 34636
rect 12597 34602 12619 34636
rect 12619 34602 12631 34636
rect 12669 34602 12687 34636
rect 12687 34602 12703 34636
rect 12741 34602 12755 34636
rect 12755 34602 12775 34636
rect 12813 34602 12823 34636
rect 12823 34602 12847 34636
rect 12885 34602 12891 34636
rect 12891 34602 12919 34636
rect 12957 34602 12959 34636
rect 12959 34602 12991 34636
rect 13029 34602 13061 34636
rect 13061 34602 13063 34636
rect 13101 34602 13129 34636
rect 13129 34602 13135 34636
rect 13173 34602 13197 34636
rect 13197 34602 13207 34636
rect 13245 34602 13265 34636
rect 13265 34602 13279 34636
rect 13317 34602 13333 34636
rect 13333 34602 13351 34636
rect 13389 34602 13401 34636
rect 13401 34602 13423 34636
rect 13461 34602 13469 34636
rect 13469 34602 13495 34636
rect 13533 34602 13537 34636
rect 13537 34602 13567 34636
rect 13605 34602 13639 34636
rect 1221 34452 1255 34474
rect 1221 34440 1255 34452
rect 1221 34384 1255 34402
rect 1221 34368 1255 34384
rect 1221 34316 1255 34330
rect 1221 34296 1255 34316
rect 1221 34248 1255 34258
rect 1221 34224 1255 34248
rect 1221 34180 1255 34186
rect 1221 34152 1255 34180
rect 1221 34112 1255 34114
rect 1221 34080 1255 34112
rect 1221 34010 1255 34042
rect 1221 34008 1255 34010
rect 1221 33942 1255 33970
rect 1221 33936 1255 33942
rect 1221 33874 1255 33898
rect 1221 33864 1255 33874
rect 1221 33806 1255 33826
rect 1221 33792 1255 33806
rect 1221 33738 1255 33754
rect 1221 33720 1255 33738
rect 1221 33670 1255 33682
rect 1221 33648 1255 33670
rect 1221 33602 1255 33610
rect 1221 33576 1255 33602
rect 1221 33534 1255 33538
rect 1221 33504 1255 33534
rect 1221 33432 1255 33466
rect 1221 33364 1255 33394
rect 1221 33360 1255 33364
rect 1221 33296 1255 33322
rect 1221 33288 1255 33296
rect 1221 33228 1255 33250
rect 1221 33216 1255 33228
rect 1221 33160 1255 33178
rect 1221 33144 1255 33160
rect 1221 33092 1255 33106
rect 1221 33072 1255 33092
rect 1221 33024 1255 33034
rect 1221 33000 1255 33024
rect 1221 32956 1255 32962
rect 1221 32928 1255 32956
rect 1221 32888 1255 32890
rect 1221 32856 1255 32888
rect 1221 32786 1255 32818
rect 1221 32784 1255 32786
rect 1221 32718 1255 32746
rect 1221 32712 1255 32718
rect 1221 32650 1255 32674
rect 1221 32640 1255 32650
rect 1221 32582 1255 32602
rect 1221 32568 1255 32582
rect 1221 32514 1255 32530
rect 1221 32496 1255 32514
rect 1221 32446 1255 32458
rect 1221 32424 1255 32446
rect 1221 32378 1255 32386
rect 1221 32352 1255 32378
rect 1221 32310 1255 32314
rect 1221 32280 1255 32310
rect 1221 32208 1255 32242
rect 1221 32140 1255 32170
rect 1221 32136 1255 32140
rect 1221 32072 1255 32098
rect 1221 32064 1255 32072
rect 1221 32004 1255 32026
rect 1221 31992 1255 32004
rect 1221 31936 1255 31954
rect 1221 31920 1255 31936
rect 1221 31868 1255 31882
rect 1221 31848 1255 31868
rect 1221 31800 1255 31810
rect 1221 31776 1255 31800
rect 1221 31732 1255 31738
rect 1221 31704 1255 31732
rect 1221 31664 1255 31666
rect 1221 31632 1255 31664
rect 1221 31562 1255 31594
rect 1221 31560 1255 31562
rect 1221 31494 1255 31522
rect 1221 31488 1255 31494
rect 1221 31426 1255 31450
rect 1221 31416 1255 31426
rect 1221 31358 1255 31378
rect 1221 31344 1255 31358
rect 1221 31290 1255 31306
rect 1221 31272 1255 31290
rect 1221 31222 1255 31234
rect 1221 31200 1255 31222
rect 1221 31154 1255 31162
rect 1221 31128 1255 31154
rect 1221 31086 1255 31090
rect 1221 31056 1255 31086
rect 1221 30984 1255 31018
rect 1221 30916 1255 30946
rect 1221 30912 1255 30916
rect 1221 30848 1255 30874
rect 1221 30840 1255 30848
rect 1221 30780 1255 30802
rect 1221 30768 1255 30780
rect 1221 30712 1255 30730
rect 1221 30696 1255 30712
rect 1221 30644 1255 30658
rect 1221 30624 1255 30644
rect 1221 30576 1255 30586
rect 1221 30552 1255 30576
rect 1221 30508 1255 30514
rect 1221 30480 1255 30508
rect 1221 30440 1255 30442
rect 1221 30408 1255 30440
rect 1221 30338 1255 30370
rect 1221 30336 1255 30338
rect 1221 30270 1255 30298
rect 1221 30264 1255 30270
rect 1221 30202 1255 30226
rect 1221 30192 1255 30202
rect 1221 30134 1255 30154
rect 1221 30120 1255 30134
rect 1221 30066 1255 30082
rect 1221 30048 1255 30066
rect 1221 29998 1255 30010
rect 1221 29976 1255 29998
rect 1221 29930 1255 29938
rect 1221 29904 1255 29930
rect 1221 29862 1255 29866
rect 1221 29832 1255 29862
rect 1221 29760 1255 29794
rect 1221 29692 1255 29722
rect 1221 29688 1255 29692
rect 1221 29624 1255 29650
rect 1221 29616 1255 29624
rect 1221 29556 1255 29578
rect 1221 29544 1255 29556
rect 1221 29488 1255 29506
rect 1221 29472 1255 29488
rect 1221 29420 1255 29434
rect 1221 29400 1255 29420
rect 1221 29352 1255 29362
rect 1221 29328 1255 29352
rect 1221 29284 1255 29290
rect 1221 29256 1255 29284
rect 1221 29216 1255 29218
rect 1221 29184 1255 29216
rect 1221 29114 1255 29146
rect 1221 29112 1255 29114
rect 1221 29046 1255 29074
rect 1221 29040 1255 29046
rect 1221 28978 1255 29002
rect 1221 28968 1255 28978
rect 1221 28910 1255 28930
rect 1221 28896 1255 28910
rect 1221 28842 1255 28858
rect 1221 28824 1255 28842
rect 1221 28774 1255 28786
rect 1221 28752 1255 28774
rect 1221 28706 1255 28714
rect 1221 28680 1255 28706
rect 1221 28638 1255 28642
rect 1221 28608 1255 28638
rect 1221 28536 1255 28570
rect 1221 28468 1255 28498
rect 1221 28464 1255 28468
rect 1221 28400 1255 28426
rect 1221 28392 1255 28400
rect 1221 28332 1255 28354
rect 1221 28320 1255 28332
rect 1221 28264 1255 28282
rect 1221 28248 1255 28264
rect 1221 28196 1255 28210
rect 1221 28176 1255 28196
rect 1221 28128 1255 28138
rect 1221 28104 1255 28128
rect 1221 28060 1255 28066
rect 1221 28032 1255 28060
rect 1221 27992 1255 27994
rect 1221 27960 1255 27992
rect 1221 27890 1255 27922
rect 1221 27888 1255 27890
rect 1221 27822 1255 27850
rect 1221 27816 1255 27822
rect 1221 27754 1255 27778
rect 1221 27744 1255 27754
rect 1221 27686 1255 27706
rect 1221 27672 1255 27686
rect 1221 27618 1255 27634
rect 1221 27600 1255 27618
rect 1221 27550 1255 27562
rect 1221 27528 1255 27550
rect 1221 27482 1255 27490
rect 1221 27456 1255 27482
rect 1221 27414 1255 27418
rect 1221 27384 1255 27414
rect 1221 27312 1255 27346
rect 1221 27244 1255 27274
rect 1221 27240 1255 27244
rect 1221 27176 1255 27202
rect 1221 27168 1255 27176
rect 1221 27108 1255 27130
rect 1221 27096 1255 27108
rect 1221 27040 1255 27058
rect 1221 27024 1255 27040
rect 1221 26972 1255 26986
rect 1221 26952 1255 26972
rect 1221 26904 1255 26914
rect 1221 26880 1255 26904
rect 1221 26836 1255 26842
rect 1221 26808 1255 26836
rect 1221 26768 1255 26770
rect 1221 26736 1255 26768
rect 1221 26666 1255 26698
rect 1221 26664 1255 26666
rect 1221 26598 1255 26626
rect 1221 26592 1255 26598
rect 1221 26530 1255 26554
rect 1221 26520 1255 26530
rect 1221 26462 1255 26482
rect 1221 26448 1255 26462
rect 1221 26394 1255 26410
rect 1221 26376 1255 26394
rect 1221 26326 1255 26338
rect 1221 26304 1255 26326
rect 1221 26258 1255 26266
rect 1221 26232 1255 26258
rect 1221 26190 1255 26194
rect 1221 26160 1255 26190
rect 1221 26088 1255 26122
rect 1221 26020 1255 26050
rect 1221 26016 1255 26020
rect 1221 25952 1255 25978
rect 1221 25944 1255 25952
rect 1221 25884 1255 25906
rect 1221 25872 1255 25884
rect 1221 25816 1255 25834
rect 1221 25800 1255 25816
rect 1221 25748 1255 25762
rect 1221 25728 1255 25748
rect 1221 25680 1255 25690
rect 1221 25656 1255 25680
rect 1221 25612 1255 25618
rect 1221 25584 1255 25612
rect 1221 25544 1255 25546
rect 1221 25512 1255 25544
rect 1221 25442 1255 25474
rect 1221 25440 1255 25442
rect 1221 25374 1255 25402
rect 1221 25368 1255 25374
rect 1221 25306 1255 25330
rect 1221 25296 1255 25306
rect 1221 25238 1255 25258
rect 1221 25224 1255 25238
rect 1221 25170 1255 25186
rect 1221 25152 1255 25170
rect 1221 25102 1255 25114
rect 1221 25080 1255 25102
rect 1221 25034 1255 25042
rect 1221 25008 1255 25034
rect 1221 24966 1255 24970
rect 1221 24936 1255 24966
rect 1221 24864 1255 24898
rect 1221 24796 1255 24826
rect 1221 24792 1255 24796
rect 1221 24728 1255 24754
rect 1221 24720 1255 24728
rect 1221 24660 1255 24682
rect 1221 24648 1255 24660
rect 1221 24592 1255 24610
rect 1221 24576 1255 24592
rect 1221 24524 1255 24538
rect 1221 24504 1255 24524
rect 1221 24456 1255 24466
rect 1221 24432 1255 24456
rect 1221 24388 1255 24394
rect 1221 24360 1255 24388
rect 1221 24320 1255 24322
rect 1221 24288 1255 24320
rect 1221 24218 1255 24250
rect 1221 24216 1255 24218
rect 1221 24150 1255 24178
rect 1221 24144 1255 24150
rect 1221 24082 1255 24106
rect 1221 24072 1255 24082
rect 1221 24014 1255 24034
rect 1221 24000 1255 24014
rect 1221 23946 1255 23962
rect 1221 23928 1255 23946
rect 1221 23878 1255 23890
rect 1221 23856 1255 23878
rect 1221 23810 1255 23818
rect 1221 23784 1255 23810
rect 1221 23742 1255 23746
rect 1221 23712 1255 23742
rect 1221 23640 1255 23674
rect 1221 23572 1255 23602
rect 1221 23568 1255 23572
rect 1221 23504 1255 23530
rect 1221 23496 1255 23504
rect 1221 23436 1255 23458
rect 1221 23424 1255 23436
rect 1221 23368 1255 23386
rect 1221 23352 1255 23368
rect 1221 23300 1255 23314
rect 1221 23280 1255 23300
rect 1221 23232 1255 23242
rect 1221 23208 1255 23232
rect 1221 23164 1255 23170
rect 1221 23136 1255 23164
rect 1221 23096 1255 23098
rect 1221 23064 1255 23096
rect 1221 22994 1255 23026
rect 1221 22992 1255 22994
rect 1221 22926 1255 22954
rect 1221 22920 1255 22926
rect 1221 22858 1255 22882
rect 1221 22848 1255 22858
rect 1221 22790 1255 22810
rect 1221 22776 1255 22790
rect 1221 22722 1255 22738
rect 1221 22704 1255 22722
rect 1221 22654 1255 22666
rect 1221 22632 1255 22654
rect 1221 22586 1255 22594
rect 1221 22560 1255 22586
rect 1221 22518 1255 22522
rect 1221 22488 1255 22518
rect 1221 22416 1255 22450
rect 1221 22348 1255 22378
rect 1221 22344 1255 22348
rect 1221 22280 1255 22306
rect 1221 22272 1255 22280
rect 1221 22212 1255 22234
rect 1221 22200 1255 22212
rect 1221 22144 1255 22162
rect 1221 22128 1255 22144
rect 1221 22076 1255 22090
rect 1221 22056 1255 22076
rect 1221 22008 1255 22018
rect 1221 21984 1255 22008
rect 1221 21940 1255 21946
rect 1221 21912 1255 21940
rect 1221 21872 1255 21874
rect 1221 21840 1255 21872
rect 1221 21770 1255 21802
rect 1221 21768 1255 21770
rect 1221 21702 1255 21730
rect 1221 21696 1255 21702
rect 1221 21634 1255 21658
rect 1221 21624 1255 21634
rect 1221 21566 1255 21586
rect 1221 21552 1255 21566
rect 1221 21498 1255 21514
rect 1221 21480 1255 21498
rect 1221 21430 1255 21442
rect 1221 21408 1255 21430
rect 1221 21362 1255 21370
rect 1221 21336 1255 21362
rect 1221 21294 1255 21298
rect 1221 21264 1255 21294
rect 1221 21192 1255 21226
rect 1221 21124 1255 21154
rect 1221 21120 1255 21124
rect 1221 21056 1255 21082
rect 1221 21048 1255 21056
rect 1221 20988 1255 21010
rect 1221 20976 1255 20988
rect 1221 20920 1255 20938
rect 1221 20904 1255 20920
rect 1221 20852 1255 20866
rect 1221 20832 1255 20852
rect 1221 20784 1255 20794
rect 1221 20760 1255 20784
rect 1221 20716 1255 20722
rect 1221 20688 1255 20716
rect 1221 20648 1255 20650
rect 1221 20616 1255 20648
rect 1221 20546 1255 20578
rect 1221 20544 1255 20546
rect 1221 20478 1255 20506
rect 1221 20472 1255 20478
rect 1221 20410 1255 20434
rect 1221 20400 1255 20410
rect 1221 20342 1255 20362
rect 1221 20328 1255 20342
rect 1221 20274 1255 20290
rect 1221 20256 1255 20274
rect 1221 20206 1255 20218
rect 1221 20184 1255 20206
rect 1221 20138 1255 20146
rect 1221 20112 1255 20138
rect 1221 20070 1255 20074
rect 1221 20040 1255 20070
rect 1221 19968 1255 20002
rect 1221 19900 1255 19930
rect 1221 19896 1255 19900
rect 1221 19832 1255 19858
rect 1221 19824 1255 19832
rect 1221 19764 1255 19786
rect 1221 19752 1255 19764
rect 1221 19696 1255 19714
rect 1221 19680 1255 19696
rect 1221 19628 1255 19642
rect 1221 19608 1255 19628
rect 1221 19560 1255 19570
rect 1221 19536 1255 19560
rect 1221 19492 1255 19498
rect 1221 19464 1255 19492
rect 1221 19424 1255 19426
rect 1221 19392 1255 19424
rect 1221 19322 1255 19354
rect 1221 19320 1255 19322
rect 1221 19254 1255 19282
rect 1221 19248 1255 19254
rect 1221 19186 1255 19210
rect 1221 19176 1255 19186
rect 1221 19118 1255 19138
rect 1221 19104 1255 19118
rect 1221 19050 1255 19066
rect 1221 19032 1255 19050
rect 1221 18982 1255 18994
rect 1221 18960 1255 18982
rect 1221 18914 1255 18922
rect 1221 18888 1255 18914
rect 1221 18846 1255 18850
rect 1221 18816 1255 18846
rect 1221 18744 1255 18778
rect 1221 18676 1255 18706
rect 1221 18672 1255 18676
rect 1221 18608 1255 18634
rect 1221 18600 1255 18608
rect 1221 18540 1255 18562
rect 1221 18528 1255 18540
rect 1221 18472 1255 18490
rect 1221 18456 1255 18472
rect 1221 18404 1255 18418
rect 1221 18384 1255 18404
rect 1221 18336 1255 18346
rect 1221 18312 1255 18336
rect 1221 18268 1255 18274
rect 1221 18240 1255 18268
rect 1221 18200 1255 18202
rect 1221 18168 1255 18200
rect 1221 18098 1255 18130
rect 1221 18096 1255 18098
rect 1221 18030 1255 18058
rect 1221 18024 1255 18030
rect 1221 17962 1255 17986
rect 1221 17952 1255 17962
rect 1221 17894 1255 17914
rect 1221 17880 1255 17894
rect 1221 17826 1255 17842
rect 1221 17808 1255 17826
rect 1221 17758 1255 17770
rect 1221 17736 1255 17758
rect 1221 17690 1255 17698
rect 1221 17664 1255 17690
rect 1221 17622 1255 17626
rect 1221 17592 1255 17622
rect 1221 17520 1255 17554
rect 1221 17452 1255 17482
rect 1221 17448 1255 17452
rect 1221 17384 1255 17410
rect 1221 17376 1255 17384
rect 1221 17316 1255 17338
rect 1221 17304 1255 17316
rect 1221 17248 1255 17266
rect 1221 17232 1255 17248
rect 1221 17180 1255 17194
rect 1221 17160 1255 17180
rect 1221 17112 1255 17122
rect 1221 17088 1255 17112
rect 1221 17044 1255 17050
rect 1221 17016 1255 17044
rect 1221 16976 1255 16978
rect 1221 16944 1255 16976
rect 1221 16874 1255 16906
rect 1221 16872 1255 16874
rect 1221 16806 1255 16834
rect 1221 16800 1255 16806
rect 1221 16738 1255 16762
rect 1221 16728 1255 16738
rect 1221 16670 1255 16690
rect 1221 16656 1255 16670
rect 1221 16602 1255 16618
rect 1221 16584 1255 16602
rect 1221 16534 1255 16546
rect 1221 16512 1255 16534
rect 1221 16466 1255 16474
rect 1221 16440 1255 16466
rect 1221 16398 1255 16402
rect 1221 16368 1255 16398
rect 1221 16296 1255 16330
rect 1221 16228 1255 16258
rect 1221 16224 1255 16228
rect 1221 16160 1255 16186
rect 1221 16152 1255 16160
rect 1221 16092 1255 16114
rect 1221 16080 1255 16092
rect 1221 16024 1255 16042
rect 1221 16008 1255 16024
rect 1221 15956 1255 15970
rect 1221 15936 1255 15956
rect 1221 15888 1255 15898
rect 1221 15864 1255 15888
rect 1221 15820 1255 15826
rect 1221 15792 1255 15820
rect 1221 15752 1255 15754
rect 1221 15720 1255 15752
rect 1221 15650 1255 15682
rect 1221 15648 1255 15650
rect 1221 15582 1255 15610
rect 1221 15576 1255 15582
rect 1221 15514 1255 15538
rect 1221 15504 1255 15514
rect 1221 15446 1255 15466
rect 1221 15432 1255 15446
rect 1221 15378 1255 15394
rect 1221 15360 1255 15378
rect 1221 15310 1255 15322
rect 1221 15288 1255 15310
rect 1221 15242 1255 15250
rect 1221 15216 1255 15242
rect 1221 15174 1255 15178
rect 1221 15144 1255 15174
rect 1221 15072 1255 15106
rect 1221 15004 1255 15034
rect 1221 15000 1255 15004
rect 1221 14936 1255 14962
rect 1221 14928 1255 14936
rect 1221 14868 1255 14890
rect 1221 14856 1255 14868
rect 1221 14800 1255 14818
rect 1221 14784 1255 14800
rect 1221 14732 1255 14746
rect 1221 14712 1255 14732
rect 1221 14664 1255 14674
rect 1221 14640 1255 14664
rect 1221 14596 1255 14602
rect 1221 14568 1255 14596
rect 1221 14528 1255 14530
rect 1221 14496 1255 14528
rect 1221 14426 1255 14458
rect 1221 14424 1255 14426
rect 1221 14358 1255 14386
rect 1221 14352 1255 14358
rect 1221 14290 1255 14314
rect 1221 14280 1255 14290
rect 1221 14222 1255 14242
rect 1221 14208 1255 14222
rect 1221 14154 1255 14170
rect 1221 14136 1255 14154
rect 1221 14086 1255 14098
rect 1221 14064 1255 14086
rect 1221 14018 1255 14026
rect 1221 13992 1255 14018
rect 1221 13950 1255 13954
rect 1221 13920 1255 13950
rect 1221 13848 1255 13882
rect 1221 13780 1255 13810
rect 1221 13776 1255 13780
rect 1221 13712 1255 13738
rect 1221 13704 1255 13712
rect 1221 13644 1255 13666
rect 1221 13632 1255 13644
rect 1221 13576 1255 13594
rect 1221 13560 1255 13576
rect 1221 13508 1255 13522
rect 1221 13488 1255 13508
rect 1221 13440 1255 13450
rect 1221 13416 1255 13440
rect 1221 13372 1255 13378
rect 1221 13344 1255 13372
rect 1221 13304 1255 13306
rect 1221 13272 1255 13304
rect 1221 13202 1255 13234
rect 1221 13200 1255 13202
rect 1221 13134 1255 13162
rect 1221 13128 1255 13134
rect 1221 13066 1255 13090
rect 1221 13056 1255 13066
rect 1221 12998 1255 13018
rect 1221 12984 1255 12998
rect 1221 12930 1255 12946
rect 1221 12912 1255 12930
rect 1221 12862 1255 12874
rect 1221 12840 1255 12862
rect 1221 12794 1255 12802
rect 1221 12768 1255 12794
rect 1221 12726 1255 12730
rect 1221 12696 1255 12726
rect 1221 12624 1255 12658
rect 1221 12556 1255 12586
rect 1221 12552 1255 12556
rect 1221 12488 1255 12514
rect 1221 12480 1255 12488
rect 1221 12420 1255 12442
rect 1221 12408 1255 12420
rect 1221 12352 1255 12370
rect 1221 12336 1255 12352
rect 1221 12284 1255 12298
rect 1221 12264 1255 12284
rect 1221 12216 1255 12226
rect 1221 12192 1255 12216
rect 1221 12148 1255 12154
rect 1221 12120 1255 12148
rect 1221 12080 1255 12082
rect 1221 12048 1255 12080
rect 1221 11978 1255 12010
rect 1221 11976 1255 11978
rect 1221 11910 1255 11938
rect 1221 11904 1255 11910
rect 1221 11842 1255 11866
rect 1221 11832 1255 11842
rect 1221 11774 1255 11794
rect 1221 11760 1255 11774
rect 1221 11706 1255 11722
rect 1221 11688 1255 11706
rect 1221 11638 1255 11650
rect 1221 11616 1255 11638
rect 1221 11570 1255 11578
rect 1221 11544 1255 11570
rect 1221 11502 1255 11506
rect 1221 11472 1255 11502
rect 1221 11400 1255 11434
rect 1221 11332 1255 11362
rect 1221 11328 1255 11332
rect 1221 11264 1255 11290
rect 1221 11256 1255 11264
rect 1221 11196 1255 11218
rect 1221 11184 1255 11196
rect 1221 11128 1255 11146
rect 1221 11112 1255 11128
rect 1221 11060 1255 11074
rect 1221 11040 1255 11060
rect 1221 10992 1255 11002
rect 1221 10968 1255 10992
rect 1221 10924 1255 10930
rect 1221 10896 1255 10924
rect 1221 10856 1255 10858
rect 1221 10824 1255 10856
rect 1221 10754 1255 10786
rect 1221 10752 1255 10754
rect 1221 10686 1255 10714
rect 1221 10680 1255 10686
rect 1221 10618 1255 10642
rect 1221 10608 1255 10618
rect 1221 10550 1255 10570
rect 1221 10536 1255 10550
rect 1221 10482 1255 10498
rect 1221 10464 1255 10482
rect 1221 10414 1255 10426
rect 1221 10392 1255 10414
rect 13739 34456 13773 34478
rect 13739 34444 13773 34456
rect 13739 34388 13773 34406
rect 13739 34372 13773 34388
rect 13739 34320 13773 34334
rect 13739 34300 13773 34320
rect 13739 34252 13773 34262
rect 13739 34228 13773 34252
rect 13739 34184 13773 34190
rect 13739 34156 13773 34184
rect 13739 34116 13773 34118
rect 13739 34084 13773 34116
rect 13739 34014 13773 34046
rect 13739 34012 13773 34014
rect 13739 33946 13773 33974
rect 13739 33940 13773 33946
rect 13739 33878 13773 33902
rect 13739 33868 13773 33878
rect 13739 33810 13773 33830
rect 13739 33796 13773 33810
rect 13739 33742 13773 33758
rect 13739 33724 13773 33742
rect 13739 33674 13773 33686
rect 13739 33652 13773 33674
rect 13739 33606 13773 33614
rect 13739 33580 13773 33606
rect 13739 33538 13773 33542
rect 13739 33508 13773 33538
rect 13739 33436 13773 33470
rect 13739 33368 13773 33398
rect 13739 33364 13773 33368
rect 13739 33300 13773 33326
rect 13739 33292 13773 33300
rect 13739 33232 13773 33254
rect 13739 33220 13773 33232
rect 13739 33164 13773 33182
rect 13739 33148 13773 33164
rect 13739 33096 13773 33110
rect 13739 33076 13773 33096
rect 13739 33028 13773 33038
rect 13739 33004 13773 33028
rect 13739 32960 13773 32966
rect 13739 32932 13773 32960
rect 13739 32892 13773 32894
rect 13739 32860 13773 32892
rect 13739 32790 13773 32822
rect 13739 32788 13773 32790
rect 13739 32722 13773 32750
rect 13739 32716 13773 32722
rect 13739 32654 13773 32678
rect 13739 32644 13773 32654
rect 13739 32586 13773 32606
rect 13739 32572 13773 32586
rect 13739 32518 13773 32534
rect 13739 32500 13773 32518
rect 13739 32450 13773 32462
rect 13739 32428 13773 32450
rect 13739 32382 13773 32390
rect 13739 32356 13773 32382
rect 13739 32314 13773 32318
rect 13739 32284 13773 32314
rect 13739 32212 13773 32246
rect 13739 32144 13773 32174
rect 13739 32140 13773 32144
rect 13739 32076 13773 32102
rect 13739 32068 13773 32076
rect 13739 32008 13773 32030
rect 13739 31996 13773 32008
rect 13739 31940 13773 31958
rect 13739 31924 13773 31940
rect 13739 31872 13773 31886
rect 13739 31852 13773 31872
rect 13739 31804 13773 31814
rect 13739 31780 13773 31804
rect 13739 31736 13773 31742
rect 13739 31708 13773 31736
rect 13739 31668 13773 31670
rect 13739 31636 13773 31668
rect 13739 31566 13773 31598
rect 13739 31564 13773 31566
rect 13739 31498 13773 31526
rect 13739 31492 13773 31498
rect 13739 31430 13773 31454
rect 13739 31420 13773 31430
rect 13739 31362 13773 31382
rect 13739 31348 13773 31362
rect 13739 31294 13773 31310
rect 13739 31276 13773 31294
rect 13739 31226 13773 31238
rect 13739 31204 13773 31226
rect 13739 31158 13773 31166
rect 13739 31132 13773 31158
rect 13739 31090 13773 31094
rect 13739 31060 13773 31090
rect 13739 30988 13773 31022
rect 13739 30920 13773 30950
rect 13739 30916 13773 30920
rect 13739 30852 13773 30878
rect 13739 30844 13773 30852
rect 13739 30784 13773 30806
rect 13739 30772 13773 30784
rect 13739 30716 13773 30734
rect 13739 30700 13773 30716
rect 13739 30648 13773 30662
rect 13739 30628 13773 30648
rect 13739 30580 13773 30590
rect 13739 30556 13773 30580
rect 13739 30512 13773 30518
rect 13739 30484 13773 30512
rect 13739 30444 13773 30446
rect 13739 30412 13773 30444
rect 13739 30342 13773 30374
rect 13739 30340 13773 30342
rect 13739 30274 13773 30302
rect 13739 30268 13773 30274
rect 13739 30206 13773 30230
rect 13739 30196 13773 30206
rect 13739 30138 13773 30158
rect 13739 30124 13773 30138
rect 13739 30070 13773 30086
rect 13739 30052 13773 30070
rect 13739 30002 13773 30014
rect 13739 29980 13773 30002
rect 13739 29934 13773 29942
rect 13739 29908 13773 29934
rect 13739 29866 13773 29870
rect 13739 29836 13773 29866
rect 13739 29764 13773 29798
rect 13739 29696 13773 29726
rect 13739 29692 13773 29696
rect 13739 29628 13773 29654
rect 13739 29620 13773 29628
rect 13739 29560 13773 29582
rect 13739 29548 13773 29560
rect 13739 29492 13773 29510
rect 13739 29476 13773 29492
rect 13739 29424 13773 29438
rect 13739 29404 13773 29424
rect 13739 29356 13773 29366
rect 13739 29332 13773 29356
rect 13739 29288 13773 29294
rect 13739 29260 13773 29288
rect 13739 29220 13773 29222
rect 13739 29188 13773 29220
rect 13739 29118 13773 29150
rect 13739 29116 13773 29118
rect 13739 29050 13773 29078
rect 13739 29044 13773 29050
rect 13739 28982 13773 29006
rect 13739 28972 13773 28982
rect 13739 28914 13773 28934
rect 13739 28900 13773 28914
rect 13739 28846 13773 28862
rect 13739 28828 13773 28846
rect 13739 28778 13773 28790
rect 13739 28756 13773 28778
rect 13739 28710 13773 28718
rect 13739 28684 13773 28710
rect 13739 28642 13773 28646
rect 13739 28612 13773 28642
rect 13739 28540 13773 28574
rect 13739 28472 13773 28502
rect 13739 28468 13773 28472
rect 13739 28404 13773 28430
rect 13739 28396 13773 28404
rect 13739 28336 13773 28358
rect 13739 28324 13773 28336
rect 13739 28268 13773 28286
rect 13739 28252 13773 28268
rect 13739 28200 13773 28214
rect 13739 28180 13773 28200
rect 13739 28132 13773 28142
rect 13739 28108 13773 28132
rect 13739 28064 13773 28070
rect 13739 28036 13773 28064
rect 13739 27996 13773 27998
rect 13739 27964 13773 27996
rect 13739 27894 13773 27926
rect 13739 27892 13773 27894
rect 13739 27826 13773 27854
rect 13739 27820 13773 27826
rect 13739 27758 13773 27782
rect 13739 27748 13773 27758
rect 13739 27690 13773 27710
rect 13739 27676 13773 27690
rect 13739 27622 13773 27638
rect 13739 27604 13773 27622
rect 13739 27554 13773 27566
rect 13739 27532 13773 27554
rect 13739 27486 13773 27494
rect 13739 27460 13773 27486
rect 13739 27418 13773 27422
rect 13739 27388 13773 27418
rect 13739 27316 13773 27350
rect 13739 27248 13773 27278
rect 13739 27244 13773 27248
rect 13739 27180 13773 27206
rect 13739 27172 13773 27180
rect 13739 27112 13773 27134
rect 13739 27100 13773 27112
rect 13739 27044 13773 27062
rect 13739 27028 13773 27044
rect 13739 26976 13773 26990
rect 13739 26956 13773 26976
rect 13739 26908 13773 26918
rect 13739 26884 13773 26908
rect 13739 26840 13773 26846
rect 13739 26812 13773 26840
rect 13739 26772 13773 26774
rect 13739 26740 13773 26772
rect 13739 26670 13773 26702
rect 13739 26668 13773 26670
rect 13739 26602 13773 26630
rect 13739 26596 13773 26602
rect 13739 26534 13773 26558
rect 13739 26524 13773 26534
rect 13739 26466 13773 26486
rect 13739 26452 13773 26466
rect 13739 26398 13773 26414
rect 13739 26380 13773 26398
rect 13739 26330 13773 26342
rect 13739 26308 13773 26330
rect 13739 26262 13773 26270
rect 13739 26236 13773 26262
rect 13739 26194 13773 26198
rect 13739 26164 13773 26194
rect 13739 26092 13773 26126
rect 13739 26024 13773 26054
rect 13739 26020 13773 26024
rect 13739 25956 13773 25982
rect 13739 25948 13773 25956
rect 13739 25888 13773 25910
rect 13739 25876 13773 25888
rect 13739 25820 13773 25838
rect 13739 25804 13773 25820
rect 13739 25752 13773 25766
rect 13739 25732 13773 25752
rect 13739 25684 13773 25694
rect 13739 25660 13773 25684
rect 13739 25616 13773 25622
rect 13739 25588 13773 25616
rect 13739 25548 13773 25550
rect 13739 25516 13773 25548
rect 13739 25446 13773 25478
rect 13739 25444 13773 25446
rect 13739 25378 13773 25406
rect 13739 25372 13773 25378
rect 13739 25310 13773 25334
rect 13739 25300 13773 25310
rect 13739 25242 13773 25262
rect 13739 25228 13773 25242
rect 13739 25174 13773 25190
rect 13739 25156 13773 25174
rect 13739 25106 13773 25118
rect 13739 25084 13773 25106
rect 13739 25038 13773 25046
rect 13739 25012 13773 25038
rect 13739 24970 13773 24974
rect 13739 24940 13773 24970
rect 13739 24868 13773 24902
rect 13739 24800 13773 24830
rect 13739 24796 13773 24800
rect 13739 24732 13773 24758
rect 13739 24724 13773 24732
rect 13739 24664 13773 24686
rect 13739 24652 13773 24664
rect 13739 24596 13773 24614
rect 13739 24580 13773 24596
rect 13739 24528 13773 24542
rect 13739 24508 13773 24528
rect 13739 24460 13773 24470
rect 13739 24436 13773 24460
rect 13739 24392 13773 24398
rect 13739 24364 13773 24392
rect 13739 24324 13773 24326
rect 13739 24292 13773 24324
rect 13739 24222 13773 24254
rect 13739 24220 13773 24222
rect 13739 24154 13773 24182
rect 13739 24148 13773 24154
rect 13739 24086 13773 24110
rect 13739 24076 13773 24086
rect 13739 24018 13773 24038
rect 13739 24004 13773 24018
rect 13739 23950 13773 23966
rect 13739 23932 13773 23950
rect 13739 23882 13773 23894
rect 13739 23860 13773 23882
rect 13739 23814 13773 23822
rect 13739 23788 13773 23814
rect 13739 23746 13773 23750
rect 13739 23716 13773 23746
rect 13739 23644 13773 23678
rect 13739 23576 13773 23606
rect 13739 23572 13773 23576
rect 13739 23508 13773 23534
rect 13739 23500 13773 23508
rect 13739 23440 13773 23462
rect 13739 23428 13773 23440
rect 13739 23372 13773 23390
rect 13739 23356 13773 23372
rect 13739 23304 13773 23318
rect 13739 23284 13773 23304
rect 13739 23236 13773 23246
rect 13739 23212 13773 23236
rect 13739 23168 13773 23174
rect 13739 23140 13773 23168
rect 13739 23100 13773 23102
rect 13739 23068 13773 23100
rect 13739 22998 13773 23030
rect 13739 22996 13773 22998
rect 13739 22930 13773 22958
rect 13739 22924 13773 22930
rect 13739 22862 13773 22886
rect 13739 22852 13773 22862
rect 13739 22794 13773 22814
rect 13739 22780 13773 22794
rect 13739 22726 13773 22742
rect 13739 22708 13773 22726
rect 13739 22658 13773 22670
rect 13739 22636 13773 22658
rect 13739 22590 13773 22598
rect 13739 22564 13773 22590
rect 13739 22522 13773 22526
rect 13739 22492 13773 22522
rect 13739 22420 13773 22454
rect 13739 22352 13773 22382
rect 13739 22348 13773 22352
rect 13739 22284 13773 22310
rect 13739 22276 13773 22284
rect 13739 22216 13773 22238
rect 13739 22204 13773 22216
rect 13739 22148 13773 22166
rect 13739 22132 13773 22148
rect 13739 22080 13773 22094
rect 13739 22060 13773 22080
rect 13739 22012 13773 22022
rect 13739 21988 13773 22012
rect 13739 21944 13773 21950
rect 13739 21916 13773 21944
rect 13739 21876 13773 21878
rect 13739 21844 13773 21876
rect 13739 21774 13773 21806
rect 13739 21772 13773 21774
rect 13739 21706 13773 21734
rect 13739 21700 13773 21706
rect 13739 21638 13773 21662
rect 13739 21628 13773 21638
rect 13739 21570 13773 21590
rect 13739 21556 13773 21570
rect 13739 21502 13773 21518
rect 13739 21484 13773 21502
rect 13739 21434 13773 21446
rect 13739 21412 13773 21434
rect 13739 21366 13773 21374
rect 13739 21340 13773 21366
rect 13739 21298 13773 21302
rect 13739 21268 13773 21298
rect 13739 21196 13773 21230
rect 13739 21128 13773 21158
rect 13739 21124 13773 21128
rect 13739 21060 13773 21086
rect 13739 21052 13773 21060
rect 13739 20992 13773 21014
rect 13739 20980 13773 20992
rect 13739 20924 13773 20942
rect 13739 20908 13773 20924
rect 13739 20856 13773 20870
rect 13739 20836 13773 20856
rect 13739 20788 13773 20798
rect 13739 20764 13773 20788
rect 13739 20720 13773 20726
rect 13739 20692 13773 20720
rect 13739 20652 13773 20654
rect 13739 20620 13773 20652
rect 13739 20550 13773 20582
rect 13739 20548 13773 20550
rect 13739 20482 13773 20510
rect 13739 20476 13773 20482
rect 13739 20414 13773 20438
rect 13739 20404 13773 20414
rect 13739 20346 13773 20366
rect 13739 20332 13773 20346
rect 13739 20278 13773 20294
rect 13739 20260 13773 20278
rect 13739 20210 13773 20222
rect 13739 20188 13773 20210
rect 13739 20142 13773 20150
rect 13739 20116 13773 20142
rect 13739 20074 13773 20078
rect 13739 20044 13773 20074
rect 13739 19972 13773 20006
rect 13739 19904 13773 19934
rect 13739 19900 13773 19904
rect 13739 19836 13773 19862
rect 13739 19828 13773 19836
rect 13739 19768 13773 19790
rect 13739 19756 13773 19768
rect 13739 19700 13773 19718
rect 13739 19684 13773 19700
rect 13739 19632 13773 19646
rect 13739 19612 13773 19632
rect 13739 19564 13773 19574
rect 13739 19540 13773 19564
rect 13739 19496 13773 19502
rect 13739 19468 13773 19496
rect 13739 19428 13773 19430
rect 13739 19396 13773 19428
rect 13739 19326 13773 19358
rect 13739 19324 13773 19326
rect 13739 19258 13773 19286
rect 13739 19252 13773 19258
rect 13739 19190 13773 19214
rect 13739 19180 13773 19190
rect 13739 19122 13773 19142
rect 13739 19108 13773 19122
rect 13739 19054 13773 19070
rect 13739 19036 13773 19054
rect 13739 18986 13773 18998
rect 13739 18964 13773 18986
rect 13739 18918 13773 18926
rect 13739 18892 13773 18918
rect 13739 18850 13773 18854
rect 13739 18820 13773 18850
rect 13739 18748 13773 18782
rect 13739 18680 13773 18710
rect 13739 18676 13773 18680
rect 13739 18612 13773 18638
rect 13739 18604 13773 18612
rect 13739 18544 13773 18566
rect 13739 18532 13773 18544
rect 13739 18476 13773 18494
rect 13739 18460 13773 18476
rect 13739 18408 13773 18422
rect 13739 18388 13773 18408
rect 13739 18340 13773 18350
rect 13739 18316 13773 18340
rect 13739 18272 13773 18278
rect 13739 18244 13773 18272
rect 13739 18204 13773 18206
rect 13739 18172 13773 18204
rect 13739 18102 13773 18134
rect 13739 18100 13773 18102
rect 13739 18034 13773 18062
rect 13739 18028 13773 18034
rect 13739 17966 13773 17990
rect 13739 17956 13773 17966
rect 13739 17898 13773 17918
rect 13739 17884 13773 17898
rect 13739 17830 13773 17846
rect 13739 17812 13773 17830
rect 13739 17762 13773 17774
rect 13739 17740 13773 17762
rect 13739 17694 13773 17702
rect 13739 17668 13773 17694
rect 13739 17626 13773 17630
rect 13739 17596 13773 17626
rect 13739 17524 13773 17558
rect 13739 17456 13773 17486
rect 13739 17452 13773 17456
rect 13739 17388 13773 17414
rect 13739 17380 13773 17388
rect 13739 17320 13773 17342
rect 13739 17308 13773 17320
rect 13739 17252 13773 17270
rect 13739 17236 13773 17252
rect 13739 17184 13773 17198
rect 13739 17164 13773 17184
rect 13739 17116 13773 17126
rect 13739 17092 13773 17116
rect 13739 17048 13773 17054
rect 13739 17020 13773 17048
rect 13739 16980 13773 16982
rect 13739 16948 13773 16980
rect 13739 16878 13773 16910
rect 13739 16876 13773 16878
rect 13739 16810 13773 16838
rect 13739 16804 13773 16810
rect 13739 16742 13773 16766
rect 13739 16732 13773 16742
rect 13739 16674 13773 16694
rect 13739 16660 13773 16674
rect 13739 16606 13773 16622
rect 13739 16588 13773 16606
rect 13739 16538 13773 16550
rect 13739 16516 13773 16538
rect 13739 16470 13773 16478
rect 13739 16444 13773 16470
rect 13739 16402 13773 16406
rect 13739 16372 13773 16402
rect 13739 16300 13773 16334
rect 13739 16232 13773 16262
rect 13739 16228 13773 16232
rect 13739 16164 13773 16190
rect 13739 16156 13773 16164
rect 13739 16096 13773 16118
rect 13739 16084 13773 16096
rect 13739 16028 13773 16046
rect 13739 16012 13773 16028
rect 13739 15960 13773 15974
rect 13739 15940 13773 15960
rect 13739 15892 13773 15902
rect 13739 15868 13773 15892
rect 13739 15824 13773 15830
rect 13739 15796 13773 15824
rect 13739 15756 13773 15758
rect 13739 15724 13773 15756
rect 13739 15654 13773 15686
rect 13739 15652 13773 15654
rect 13739 15586 13773 15614
rect 13739 15580 13773 15586
rect 13739 15518 13773 15542
rect 13739 15508 13773 15518
rect 13739 15450 13773 15470
rect 13739 15436 13773 15450
rect 13739 15382 13773 15398
rect 13739 15364 13773 15382
rect 13739 15314 13773 15326
rect 13739 15292 13773 15314
rect 13739 15246 13773 15254
rect 13739 15220 13773 15246
rect 13739 15178 13773 15182
rect 13739 15148 13773 15178
rect 13739 15076 13773 15110
rect 13739 15008 13773 15038
rect 13739 15004 13773 15008
rect 13739 14940 13773 14966
rect 13739 14932 13773 14940
rect 13739 14872 13773 14894
rect 13739 14860 13773 14872
rect 13739 14804 13773 14822
rect 13739 14788 13773 14804
rect 13739 14736 13773 14750
rect 13739 14716 13773 14736
rect 13739 14668 13773 14678
rect 13739 14644 13773 14668
rect 13739 14600 13773 14606
rect 13739 14572 13773 14600
rect 13739 14532 13773 14534
rect 13739 14500 13773 14532
rect 13739 14430 13773 14462
rect 13739 14428 13773 14430
rect 13739 14362 13773 14390
rect 13739 14356 13773 14362
rect 13739 14294 13773 14318
rect 13739 14284 13773 14294
rect 13739 14226 13773 14246
rect 13739 14212 13773 14226
rect 13739 14158 13773 14174
rect 13739 14140 13773 14158
rect 13739 14090 13773 14102
rect 13739 14068 13773 14090
rect 13739 14022 13773 14030
rect 13739 13996 13773 14022
rect 13739 13954 13773 13958
rect 13739 13924 13773 13954
rect 13739 13852 13773 13886
rect 13739 13784 13773 13814
rect 13739 13780 13773 13784
rect 13739 13716 13773 13742
rect 13739 13708 13773 13716
rect 13739 13648 13773 13670
rect 13739 13636 13773 13648
rect 13739 13580 13773 13598
rect 13739 13564 13773 13580
rect 13739 13512 13773 13526
rect 13739 13492 13773 13512
rect 13739 13444 13773 13454
rect 13739 13420 13773 13444
rect 13739 13376 13773 13382
rect 13739 13348 13773 13376
rect 13739 13308 13773 13310
rect 13739 13276 13773 13308
rect 13739 13206 13773 13238
rect 13739 13204 13773 13206
rect 13739 13138 13773 13166
rect 13739 13132 13773 13138
rect 13739 13070 13773 13094
rect 13739 13060 13773 13070
rect 13739 13002 13773 13022
rect 13739 12988 13773 13002
rect 13739 12934 13773 12950
rect 13739 12916 13773 12934
rect 13739 12866 13773 12878
rect 13739 12844 13773 12866
rect 13739 12798 13773 12806
rect 13739 12772 13773 12798
rect 13739 12730 13773 12734
rect 13739 12700 13773 12730
rect 13739 12628 13773 12662
rect 13739 12560 13773 12590
rect 13739 12556 13773 12560
rect 13739 12492 13773 12518
rect 13739 12484 13773 12492
rect 13739 12424 13773 12446
rect 13739 12412 13773 12424
rect 13739 12356 13773 12374
rect 13739 12340 13773 12356
rect 13739 12288 13773 12302
rect 13739 12268 13773 12288
rect 13739 12220 13773 12230
rect 13739 12196 13773 12220
rect 13739 12152 13773 12158
rect 13739 12124 13773 12152
rect 13739 12084 13773 12086
rect 13739 12052 13773 12084
rect 13739 11982 13773 12014
rect 13739 11980 13773 11982
rect 13739 11914 13773 11942
rect 13739 11908 13773 11914
rect 13739 11846 13773 11870
rect 13739 11836 13773 11846
rect 13739 11778 13773 11798
rect 13739 11764 13773 11778
rect 13739 11710 13773 11726
rect 13739 11692 13773 11710
rect 13739 11642 13773 11654
rect 13739 11620 13773 11642
rect 13739 11574 13773 11582
rect 13739 11548 13773 11574
rect 13739 11506 13773 11510
rect 13739 11476 13773 11506
rect 13739 11404 13773 11438
rect 13739 11336 13773 11366
rect 13739 11332 13773 11336
rect 13739 11268 13773 11294
rect 13739 11260 13773 11268
rect 13739 11200 13773 11222
rect 13739 11188 13773 11200
rect 13739 11132 13773 11150
rect 13739 11116 13773 11132
rect 13739 11064 13773 11078
rect 13739 11044 13773 11064
rect 13739 10996 13773 11006
rect 13739 10972 13773 10996
rect 13739 10928 13773 10934
rect 13739 10900 13773 10928
rect 13739 10860 13773 10862
rect 13739 10828 13773 10860
rect 13739 10758 13773 10790
rect 13739 10756 13773 10758
rect 13739 10690 13773 10718
rect 13739 10684 13773 10690
rect 13739 10622 13773 10646
rect 13739 10612 13773 10622
rect 13739 10554 13773 10574
rect 13739 10540 13773 10554
rect 13739 10486 13773 10502
rect 13739 10468 13773 10486
rect 13739 10418 13773 10430
rect 13739 10396 13773 10418
rect 1355 10256 1389 10290
rect 1427 10256 1457 10290
rect 1457 10256 1461 10290
rect 1499 10256 1525 10290
rect 1525 10256 1533 10290
rect 1571 10256 1593 10290
rect 1593 10256 1605 10290
rect 1643 10256 1661 10290
rect 1661 10256 1677 10290
rect 1715 10256 1729 10290
rect 1729 10256 1749 10290
rect 1787 10256 1797 10290
rect 1797 10256 1821 10290
rect 1859 10256 1865 10290
rect 1865 10256 1893 10290
rect 1931 10256 1933 10290
rect 1933 10256 1965 10290
rect 2003 10256 2035 10290
rect 2035 10256 2037 10290
rect 2075 10256 2103 10290
rect 2103 10256 2109 10290
rect 2147 10256 2171 10290
rect 2171 10256 2181 10290
rect 2219 10256 2239 10290
rect 2239 10256 2253 10290
rect 2291 10256 2307 10290
rect 2307 10256 2325 10290
rect 2363 10256 2375 10290
rect 2375 10256 2397 10290
rect 2435 10256 2443 10290
rect 2443 10256 2469 10290
rect 2507 10256 2511 10290
rect 2511 10256 2541 10290
rect 2579 10256 2613 10290
rect 2651 10256 2681 10290
rect 2681 10256 2685 10290
rect 2723 10256 2749 10290
rect 2749 10256 2757 10290
rect 2795 10256 2817 10290
rect 2817 10256 2829 10290
rect 2867 10256 2885 10290
rect 2885 10256 2901 10290
rect 2939 10256 2953 10290
rect 2953 10256 2973 10290
rect 3011 10256 3021 10290
rect 3021 10256 3045 10290
rect 3083 10256 3089 10290
rect 3089 10256 3117 10290
rect 3155 10256 3157 10290
rect 3157 10256 3189 10290
rect 3227 10256 3259 10290
rect 3259 10256 3261 10290
rect 3299 10256 3327 10290
rect 3327 10256 3333 10290
rect 3371 10256 3395 10290
rect 3395 10256 3405 10290
rect 3443 10256 3463 10290
rect 3463 10256 3477 10290
rect 3515 10256 3531 10290
rect 3531 10256 3549 10290
rect 3587 10256 3599 10290
rect 3599 10256 3621 10290
rect 3659 10256 3667 10290
rect 3667 10256 3693 10290
rect 3731 10256 3735 10290
rect 3735 10256 3765 10290
rect 3803 10256 3837 10290
rect 3875 10256 3905 10290
rect 3905 10256 3909 10290
rect 3947 10256 3973 10290
rect 3973 10256 3981 10290
rect 4019 10256 4041 10290
rect 4041 10256 4053 10290
rect 4091 10256 4109 10290
rect 4109 10256 4125 10290
rect 4163 10256 4177 10290
rect 4177 10256 4197 10290
rect 4235 10256 4245 10290
rect 4245 10256 4269 10290
rect 4307 10256 4313 10290
rect 4313 10256 4341 10290
rect 4379 10256 4381 10290
rect 4381 10256 4413 10290
rect 4451 10256 4483 10290
rect 4483 10256 4485 10290
rect 4523 10256 4551 10290
rect 4551 10256 4557 10290
rect 4595 10256 4619 10290
rect 4619 10256 4629 10290
rect 4667 10256 4687 10290
rect 4687 10256 4701 10290
rect 4739 10256 4755 10290
rect 4755 10256 4773 10290
rect 4811 10256 4823 10290
rect 4823 10256 4845 10290
rect 4883 10256 4891 10290
rect 4891 10256 4917 10290
rect 4955 10256 4959 10290
rect 4959 10256 4989 10290
rect 5027 10256 5061 10290
rect 5099 10256 5129 10290
rect 5129 10256 5133 10290
rect 5171 10256 5197 10290
rect 5197 10256 5205 10290
rect 5243 10256 5265 10290
rect 5265 10256 5277 10290
rect 5315 10256 5333 10290
rect 5333 10256 5349 10290
rect 5387 10256 5401 10290
rect 5401 10256 5421 10290
rect 5459 10256 5469 10290
rect 5469 10256 5493 10290
rect 5531 10256 5537 10290
rect 5537 10256 5565 10290
rect 5603 10256 5605 10290
rect 5605 10256 5637 10290
rect 5675 10256 5707 10290
rect 5707 10256 5709 10290
rect 5747 10256 5775 10290
rect 5775 10256 5781 10290
rect 5819 10256 5843 10290
rect 5843 10256 5853 10290
rect 5891 10256 5911 10290
rect 5911 10256 5925 10290
rect 5963 10256 5979 10290
rect 5979 10256 5997 10290
rect 6035 10256 6047 10290
rect 6047 10256 6069 10290
rect 6107 10256 6115 10290
rect 6115 10256 6141 10290
rect 6179 10256 6183 10290
rect 6183 10256 6213 10290
rect 6251 10256 6285 10290
rect 6323 10256 6353 10290
rect 6353 10256 6357 10290
rect 6395 10256 6421 10290
rect 6421 10256 6429 10290
rect 6467 10256 6489 10290
rect 6489 10256 6501 10290
rect 6539 10256 6557 10290
rect 6557 10256 6573 10290
rect 6611 10256 6625 10290
rect 6625 10256 6645 10290
rect 6683 10256 6693 10290
rect 6693 10256 6717 10290
rect 6755 10256 6761 10290
rect 6761 10256 6789 10290
rect 6827 10256 6829 10290
rect 6829 10256 6861 10290
rect 6899 10256 6931 10290
rect 6931 10256 6933 10290
rect 6971 10256 6999 10290
rect 6999 10256 7005 10290
rect 7043 10256 7067 10290
rect 7067 10256 7077 10290
rect 7115 10256 7135 10290
rect 7135 10256 7149 10290
rect 7187 10256 7203 10290
rect 7203 10256 7221 10290
rect 7259 10256 7271 10290
rect 7271 10256 7293 10290
rect 7331 10256 7339 10290
rect 7339 10256 7365 10290
rect 7403 10256 7407 10290
rect 7407 10256 7437 10290
rect 7475 10256 7509 10290
rect 7547 10256 7577 10290
rect 7577 10256 7581 10290
rect 7619 10256 7645 10290
rect 7645 10256 7653 10290
rect 7691 10256 7713 10290
rect 7713 10256 7725 10290
rect 7763 10256 7781 10290
rect 7781 10256 7797 10290
rect 7835 10256 7849 10290
rect 7849 10256 7869 10290
rect 7907 10256 7917 10290
rect 7917 10256 7941 10290
rect 7979 10256 7985 10290
rect 7985 10256 8013 10290
rect 8051 10256 8053 10290
rect 8053 10256 8085 10290
rect 8123 10256 8155 10290
rect 8155 10256 8157 10290
rect 8195 10256 8223 10290
rect 8223 10256 8229 10290
rect 8267 10256 8291 10290
rect 8291 10256 8301 10290
rect 8339 10256 8359 10290
rect 8359 10256 8373 10290
rect 8411 10256 8427 10290
rect 8427 10256 8445 10290
rect 8483 10256 8495 10290
rect 8495 10256 8517 10290
rect 8555 10256 8563 10290
rect 8563 10256 8589 10290
rect 8627 10256 8631 10290
rect 8631 10256 8661 10290
rect 8699 10256 8733 10290
rect 8771 10256 8801 10290
rect 8801 10256 8805 10290
rect 8843 10256 8869 10290
rect 8869 10256 8877 10290
rect 8915 10256 8937 10290
rect 8937 10256 8949 10290
rect 8987 10256 9005 10290
rect 9005 10256 9021 10290
rect 9059 10256 9073 10290
rect 9073 10256 9093 10290
rect 9131 10256 9141 10290
rect 9141 10256 9165 10290
rect 9203 10256 9209 10290
rect 9209 10256 9237 10290
rect 9275 10256 9277 10290
rect 9277 10256 9309 10290
rect 9347 10256 9379 10290
rect 9379 10256 9381 10290
rect 9419 10256 9447 10290
rect 9447 10256 9453 10290
rect 9491 10256 9515 10290
rect 9515 10256 9525 10290
rect 9563 10256 9583 10290
rect 9583 10256 9597 10290
rect 9635 10256 9651 10290
rect 9651 10256 9669 10290
rect 9707 10256 9719 10290
rect 9719 10256 9741 10290
rect 9779 10256 9787 10290
rect 9787 10256 9813 10290
rect 9851 10256 9855 10290
rect 9855 10256 9885 10290
rect 9923 10256 9957 10290
rect 9995 10256 10025 10290
rect 10025 10256 10029 10290
rect 10067 10256 10093 10290
rect 10093 10256 10101 10290
rect 10139 10256 10161 10290
rect 10161 10256 10173 10290
rect 10211 10256 10229 10290
rect 10229 10256 10245 10290
rect 10283 10256 10297 10290
rect 10297 10256 10317 10290
rect 10355 10256 10365 10290
rect 10365 10256 10389 10290
rect 10427 10256 10433 10290
rect 10433 10256 10461 10290
rect 10499 10256 10501 10290
rect 10501 10256 10533 10290
rect 10571 10256 10603 10290
rect 10603 10256 10605 10290
rect 10643 10256 10671 10290
rect 10671 10256 10677 10290
rect 10715 10256 10739 10290
rect 10739 10256 10749 10290
rect 10787 10256 10807 10290
rect 10807 10256 10821 10290
rect 10859 10256 10875 10290
rect 10875 10256 10893 10290
rect 10931 10256 10943 10290
rect 10943 10256 10965 10290
rect 11003 10256 11011 10290
rect 11011 10256 11037 10290
rect 11075 10256 11079 10290
rect 11079 10256 11109 10290
rect 11147 10256 11181 10290
rect 11219 10256 11249 10290
rect 11249 10256 11253 10290
rect 11291 10256 11317 10290
rect 11317 10256 11325 10290
rect 11363 10256 11385 10290
rect 11385 10256 11397 10290
rect 11435 10256 11453 10290
rect 11453 10256 11469 10290
rect 11507 10256 11521 10290
rect 11521 10256 11541 10290
rect 11579 10256 11589 10290
rect 11589 10256 11613 10290
rect 11651 10256 11657 10290
rect 11657 10256 11685 10290
rect 11723 10256 11725 10290
rect 11725 10256 11757 10290
rect 11795 10256 11827 10290
rect 11827 10256 11829 10290
rect 11867 10256 11895 10290
rect 11895 10256 11901 10290
rect 11939 10256 11963 10290
rect 11963 10256 11973 10290
rect 12011 10256 12031 10290
rect 12031 10256 12045 10290
rect 12083 10256 12099 10290
rect 12099 10256 12117 10290
rect 12155 10256 12167 10290
rect 12167 10256 12189 10290
rect 12227 10256 12235 10290
rect 12235 10256 12261 10290
rect 12299 10256 12303 10290
rect 12303 10256 12333 10290
rect 12371 10256 12405 10290
rect 12443 10256 12473 10290
rect 12473 10256 12477 10290
rect 12515 10256 12541 10290
rect 12541 10256 12549 10290
rect 12587 10256 12609 10290
rect 12609 10256 12621 10290
rect 12659 10256 12677 10290
rect 12677 10256 12693 10290
rect 12731 10256 12745 10290
rect 12745 10256 12765 10290
rect 12803 10256 12813 10290
rect 12813 10256 12837 10290
rect 12875 10256 12881 10290
rect 12881 10256 12909 10290
rect 12947 10256 12949 10290
rect 12949 10256 12981 10290
rect 13019 10256 13051 10290
rect 13051 10256 13053 10290
rect 13091 10256 13119 10290
rect 13119 10256 13125 10290
rect 13163 10256 13187 10290
rect 13187 10256 13197 10290
rect 13235 10256 13255 10290
rect 13255 10256 13269 10290
rect 13307 10256 13323 10290
rect 13323 10256 13341 10290
rect 13379 10256 13391 10290
rect 13391 10256 13413 10290
rect 13451 10256 13459 10290
rect 13459 10256 13485 10290
rect 13523 10256 13527 10290
rect 13527 10256 13557 10290
rect 13595 10256 13629 10290
rect 14120 34646 14154 34680
rect 14120 34574 14154 34608
rect 14120 34502 14154 34536
rect 14120 34430 14154 34464
rect 14120 34358 14154 34392
rect 14120 34286 14154 34320
rect 14120 34214 14154 34248
rect 14120 34142 14154 34176
rect 14120 34070 14154 34104
rect 14120 33998 14154 34032
rect 14120 33926 14154 33960
rect 14120 33854 14154 33888
rect 14120 33782 14154 33816
rect 14120 33710 14154 33744
rect 14120 33638 14154 33672
rect 14120 33566 14154 33600
rect 14120 33494 14154 33528
rect 14120 33422 14154 33456
rect 14120 33350 14154 33384
rect 14120 33278 14154 33312
rect 14120 33206 14154 33240
rect 14120 33134 14154 33168
rect 14120 33062 14154 33096
rect 14120 32990 14154 33024
rect 14120 32918 14154 32952
rect 14120 32846 14154 32880
rect 14120 32774 14154 32808
rect 14120 32702 14154 32736
rect 14120 32630 14154 32664
rect 14120 32558 14154 32592
rect 14120 32486 14154 32520
rect 14120 32414 14154 32448
rect 14120 32342 14154 32376
rect 14120 32270 14154 32304
rect 14120 32198 14154 32232
rect 14120 32126 14154 32160
rect 14120 32054 14154 32088
rect 14120 31982 14154 32016
rect 14120 31910 14154 31944
rect 14120 31838 14154 31872
rect 14120 31766 14154 31800
rect 14120 31694 14154 31728
rect 14120 31622 14154 31656
rect 14120 31550 14154 31584
rect 14120 31478 14154 31512
rect 14120 31406 14154 31440
rect 14120 31334 14154 31368
rect 14120 31262 14154 31296
rect 14120 31190 14154 31224
rect 14120 31118 14154 31152
rect 14120 31046 14154 31080
rect 14120 30974 14154 31008
rect 14120 30902 14154 30936
rect 14120 30830 14154 30864
rect 14120 30758 14154 30792
rect 14120 30686 14154 30720
rect 14120 30614 14154 30648
rect 14120 30542 14154 30576
rect 14120 30470 14154 30504
rect 14120 30398 14154 30432
rect 14120 30326 14154 30360
rect 14120 30254 14154 30288
rect 14120 30182 14154 30216
rect 14120 30110 14154 30144
rect 14120 30038 14154 30072
rect 14120 29966 14154 30000
rect 14120 29894 14154 29928
rect 14120 29822 14154 29856
rect 14120 29750 14154 29784
rect 14120 29678 14154 29712
rect 14120 29606 14154 29640
rect 14120 29534 14154 29568
rect 14120 29462 14154 29496
rect 14120 29390 14154 29424
rect 14120 29318 14154 29352
rect 14120 29246 14154 29280
rect 14120 29174 14154 29208
rect 14120 29102 14154 29136
rect 14120 29030 14154 29064
rect 14120 28958 14154 28992
rect 14120 28886 14154 28920
rect 14120 28814 14154 28848
rect 14120 28742 14154 28776
rect 14120 28670 14154 28704
rect 14120 28598 14154 28632
rect 14120 28526 14154 28560
rect 14120 28454 14154 28488
rect 14120 28382 14154 28416
rect 14120 28310 14154 28344
rect 14120 28238 14154 28272
rect 14120 28166 14154 28200
rect 14120 28094 14154 28128
rect 14120 28022 14154 28056
rect 14120 27950 14154 27984
rect 14120 27878 14154 27912
rect 14120 27806 14154 27840
rect 14120 27734 14154 27768
rect 14120 27662 14154 27696
rect 14120 27590 14154 27624
rect 14120 27518 14154 27552
rect 14120 27446 14154 27480
rect 14120 27374 14154 27408
rect 14120 27302 14154 27336
rect 14120 27230 14154 27264
rect 14120 27158 14154 27192
rect 14120 27086 14154 27120
rect 14120 27014 14154 27048
rect 14120 26942 14154 26976
rect 14120 26870 14154 26904
rect 14120 26798 14154 26832
rect 14120 26726 14154 26760
rect 14120 26654 14154 26688
rect 14120 26582 14154 26616
rect 14120 26510 14154 26544
rect 14120 26438 14154 26472
rect 14120 26366 14154 26400
rect 14120 26294 14154 26328
rect 14120 26222 14154 26256
rect 14120 26150 14154 26184
rect 14120 26078 14154 26112
rect 14120 26006 14154 26040
rect 14120 25934 14154 25968
rect 14120 25862 14154 25896
rect 14120 25790 14154 25824
rect 14120 25718 14154 25752
rect 14120 25646 14154 25680
rect 14120 25574 14154 25608
rect 14120 25502 14154 25536
rect 14120 25430 14154 25464
rect 14120 25358 14154 25392
rect 14120 25286 14154 25320
rect 14120 25214 14154 25248
rect 14120 25142 14154 25176
rect 14120 25070 14154 25104
rect 14120 24998 14154 25032
rect 14120 24926 14154 24960
rect 14120 24854 14154 24888
rect 14120 24782 14154 24816
rect 14120 24710 14154 24744
rect 14120 24638 14154 24672
rect 14120 24566 14154 24600
rect 14120 24494 14154 24528
rect 14120 24422 14154 24456
rect 14120 24350 14154 24384
rect 14120 24278 14154 24312
rect 14120 24206 14154 24240
rect 14120 24134 14154 24168
rect 14120 24062 14154 24096
rect 14120 23990 14154 24024
rect 14120 23918 14154 23952
rect 14120 23846 14154 23880
rect 14120 23774 14154 23808
rect 14120 23702 14154 23736
rect 14120 23630 14154 23664
rect 14120 23558 14154 23592
rect 14120 23486 14154 23520
rect 14120 23414 14154 23448
rect 14120 23342 14154 23376
rect 14120 23270 14154 23304
rect 14120 23198 14154 23232
rect 14120 23126 14154 23160
rect 14120 23054 14154 23088
rect 14120 22982 14154 23016
rect 14120 22910 14154 22944
rect 14120 22838 14154 22872
rect 14120 22766 14154 22800
rect 14120 22694 14154 22728
rect 14120 22622 14154 22656
rect 14120 22550 14154 22584
rect 14120 22478 14154 22512
rect 14120 22406 14154 22440
rect 14120 22334 14154 22368
rect 14120 22262 14154 22296
rect 14120 22190 14154 22224
rect 14120 22118 14154 22152
rect 14120 22046 14154 22080
rect 14120 21974 14154 22008
rect 14120 21902 14154 21936
rect 14120 21830 14154 21864
rect 14120 21758 14154 21792
rect 14120 21686 14154 21720
rect 14120 21614 14154 21648
rect 14120 21542 14154 21576
rect 14120 21470 14154 21504
rect 14120 21398 14154 21432
rect 14120 21326 14154 21360
rect 14120 21254 14154 21288
rect 14120 21182 14154 21216
rect 14120 21110 14154 21144
rect 14120 21038 14154 21072
rect 14120 20966 14154 21000
rect 14120 20894 14154 20928
rect 14120 20822 14154 20856
rect 14120 20750 14154 20784
rect 14120 20678 14154 20712
rect 14120 20606 14154 20640
rect 14120 20534 14154 20568
rect 14120 20462 14154 20496
rect 14120 20390 14154 20424
rect 14120 20318 14154 20352
rect 14120 20246 14154 20280
rect 14120 20174 14154 20208
rect 14120 20102 14154 20136
rect 14120 20030 14154 20064
rect 14120 19958 14154 19992
rect 14120 19886 14154 19920
rect 14120 19814 14154 19848
rect 14120 19742 14154 19776
rect 14120 19670 14154 19704
rect 14120 19598 14154 19632
rect 14120 19526 14154 19560
rect 14120 19454 14154 19488
rect 14120 19382 14154 19416
rect 14120 19310 14154 19344
rect 14120 19238 14154 19272
rect 14120 19166 14154 19200
rect 14120 19094 14154 19128
rect 14120 19022 14154 19056
rect 14120 18950 14154 18984
rect 14120 18878 14154 18912
rect 14120 18806 14154 18840
rect 14120 18734 14154 18768
rect 14120 18662 14154 18696
rect 14120 18590 14154 18624
rect 14120 18518 14154 18552
rect 14120 18446 14154 18480
rect 14120 18374 14154 18408
rect 14120 18302 14154 18336
rect 14120 18230 14154 18264
rect 14120 18158 14154 18192
rect 14120 18086 14154 18120
rect 14120 18014 14154 18048
rect 14120 17942 14154 17976
rect 14120 17870 14154 17904
rect 14120 17798 14154 17832
rect 14120 17726 14154 17760
rect 14120 17654 14154 17688
rect 14120 17582 14154 17616
rect 14120 17510 14154 17544
rect 14120 17438 14154 17472
rect 14120 17366 14154 17400
rect 14120 17294 14154 17328
rect 14120 17222 14154 17256
rect 14120 17150 14154 17184
rect 14120 17078 14154 17112
rect 14120 17006 14154 17040
rect 14120 16934 14154 16968
rect 14120 16862 14154 16896
rect 14120 16790 14154 16824
rect 14120 16718 14154 16752
rect 14120 16646 14154 16680
rect 14120 16574 14154 16608
rect 14120 16502 14154 16536
rect 14120 16430 14154 16464
rect 14120 16358 14154 16392
rect 14120 16286 14154 16320
rect 14120 16214 14154 16248
rect 14120 16142 14154 16176
rect 14120 16070 14154 16104
rect 14120 15998 14154 16032
rect 14120 15926 14154 15960
rect 14120 15854 14154 15888
rect 14120 15782 14154 15816
rect 14120 15710 14154 15744
rect 14120 15638 14154 15672
rect 14120 15566 14154 15600
rect 14120 15494 14154 15528
rect 14120 15422 14154 15456
rect 14120 15350 14154 15384
rect 14120 15278 14154 15312
rect 14120 15206 14154 15240
rect 14120 15134 14154 15168
rect 14120 15062 14154 15096
rect 14120 14990 14154 15024
rect 14120 14918 14154 14952
rect 14120 14846 14154 14880
rect 14120 14774 14154 14808
rect 14120 14702 14154 14736
rect 14120 14630 14154 14664
rect 14120 14558 14154 14592
rect 14120 14486 14154 14520
rect 14120 14414 14154 14448
rect 14120 14342 14154 14376
rect 14120 14270 14154 14304
rect 14120 14198 14154 14232
rect 14120 14126 14154 14160
rect 14120 14054 14154 14088
rect 14120 13982 14154 14016
rect 14120 13910 14154 13944
rect 14120 13838 14154 13872
rect 14120 13766 14154 13800
rect 14120 13694 14154 13728
rect 14120 13622 14154 13656
rect 14120 13550 14154 13584
rect 14120 13478 14154 13512
rect 14120 13406 14154 13440
rect 14120 13334 14154 13368
rect 14120 13262 14154 13296
rect 14120 13190 14154 13224
rect 14120 13118 14154 13152
rect 14120 13046 14154 13080
rect 14120 12974 14154 13008
rect 14120 12902 14154 12936
rect 14120 12830 14154 12864
rect 14120 12758 14154 12792
rect 14120 12686 14154 12720
rect 14120 12614 14154 12648
rect 14120 12542 14154 12576
rect 14120 12470 14154 12504
rect 14120 12398 14154 12432
rect 14120 12326 14154 12360
rect 14120 12254 14154 12288
rect 14120 12182 14154 12216
rect 14120 12110 14154 12144
rect 14120 12038 14154 12072
rect 14120 11966 14154 12000
rect 14120 11894 14154 11928
rect 14120 11822 14154 11856
rect 14120 11750 14154 11784
rect 14120 11678 14154 11712
rect 14120 11606 14154 11640
rect 14120 11534 14154 11568
rect 14120 11462 14154 11496
rect 14120 11390 14154 11424
rect 14120 11318 14154 11352
rect 14120 11246 14154 11280
rect 14120 11174 14154 11208
rect 14120 11102 14154 11136
rect 14120 11030 14154 11064
rect 14120 10958 14154 10992
rect 14120 10886 14154 10920
rect 14120 10814 14154 10848
rect 14120 10742 14154 10776
rect 14120 10670 14154 10704
rect 14120 10598 14154 10632
rect 14120 10526 14154 10560
rect 14120 10454 14154 10488
rect 14120 10382 14154 10416
rect 14120 10310 14154 10344
rect 14120 10238 14154 10272
rect 814 10173 848 10207
rect 814 10101 848 10135
rect 14120 10166 14154 10200
rect 14120 10094 14154 10128
rect 912 9908 946 9942
rect 984 9908 1018 9942
rect 1056 9908 1090 9942
rect 1128 9908 1162 9942
rect 1200 9908 1234 9942
rect 1272 9908 1306 9942
rect 1344 9908 1378 9942
rect 1416 9908 1450 9942
rect 1488 9908 1522 9942
rect 1560 9908 1594 9942
rect 1632 9908 1666 9942
rect 1704 9908 1738 9942
rect 1776 9908 1810 9942
rect 1848 9908 1882 9942
rect 1920 9908 1954 9942
rect 1992 9908 2026 9942
rect 2064 9908 2098 9942
rect 2136 9908 2170 9942
rect 2208 9908 2242 9942
rect 2280 9908 2314 9942
rect 2352 9908 2386 9942
rect 2424 9908 2458 9942
rect 2496 9908 2530 9942
rect 2568 9908 2602 9942
rect 2640 9908 2674 9942
rect 2712 9908 2746 9942
rect 2784 9908 2818 9942
rect 2856 9908 2890 9942
rect 2928 9908 2962 9942
rect 3000 9908 3034 9942
rect 3072 9908 3106 9942
rect 3144 9908 3178 9942
rect 3216 9908 3250 9942
rect 3288 9908 3322 9942
rect 3360 9908 3394 9942
rect 3432 9908 3466 9942
rect 3504 9908 3538 9942
rect 3576 9908 3610 9942
rect 3648 9908 3682 9942
rect 3720 9908 3754 9942
rect 3792 9908 3826 9942
rect 3864 9908 3898 9942
rect 3936 9908 3970 9942
rect 4008 9908 4042 9942
rect 4080 9908 4114 9942
rect 4152 9908 4186 9942
rect 4224 9908 4258 9942
rect 4296 9908 4330 9942
rect 4368 9908 4402 9942
rect 4440 9908 4474 9942
rect 4512 9908 4546 9942
rect 4584 9908 4618 9942
rect 4656 9908 4690 9942
rect 4728 9908 4762 9942
rect 4800 9908 4834 9942
rect 4872 9908 4906 9942
rect 4944 9908 4978 9942
rect 5016 9908 5050 9942
rect 5088 9908 5122 9942
rect 5160 9908 5194 9942
rect 5232 9908 5266 9942
rect 5304 9908 5338 9942
rect 5376 9908 5410 9942
rect 5448 9908 5482 9942
rect 5520 9908 5554 9942
rect 5592 9908 5626 9942
rect 5664 9908 5698 9942
rect 5736 9908 5770 9942
rect 5808 9908 5842 9942
rect 5880 9908 5914 9942
rect 5952 9908 5986 9942
rect 6024 9908 6058 9942
rect 6096 9908 6130 9942
rect 6168 9908 6202 9942
rect 6240 9908 6274 9942
rect 6312 9908 6346 9942
rect 6384 9908 6418 9942
rect 6456 9908 6490 9942
rect 6528 9908 6562 9942
rect 6600 9908 6634 9942
rect 6672 9908 6706 9942
rect 6744 9908 6778 9942
rect 6816 9908 6850 9942
rect 6888 9908 6922 9942
rect 6960 9908 6994 9942
rect 7032 9908 7066 9942
rect 7104 9908 7138 9942
rect 7176 9908 7210 9942
rect 7248 9908 7282 9942
rect 7320 9908 7354 9942
rect 7392 9908 7426 9942
rect 7464 9908 7498 9942
rect 7536 9908 7570 9942
rect 7608 9908 7642 9942
rect 7680 9908 7714 9942
rect 7752 9908 7786 9942
rect 7824 9908 7858 9942
rect 7896 9908 7930 9942
rect 7968 9908 8002 9942
rect 8040 9908 8074 9942
rect 8112 9908 8146 9942
rect 8184 9908 8218 9942
rect 8256 9908 8290 9942
rect 8328 9908 8362 9942
rect 8400 9908 8434 9942
rect 8472 9908 8506 9942
rect 8544 9908 8578 9942
rect 8616 9908 8650 9942
rect 8688 9908 8722 9942
rect 8760 9908 8794 9942
rect 8832 9908 8866 9942
rect 8904 9908 8938 9942
rect 8976 9908 9010 9942
rect 9048 9908 9082 9942
rect 9120 9908 9154 9942
rect 9192 9908 9226 9942
rect 9264 9908 9298 9942
rect 9336 9908 9370 9942
rect 9408 9908 9442 9942
rect 9480 9908 9514 9942
rect 9552 9908 9586 9942
rect 9624 9908 9658 9942
rect 9696 9908 9730 9942
rect 9768 9908 9802 9942
rect 9840 9908 9874 9942
rect 9912 9908 9946 9942
rect 9984 9908 10018 9942
rect 10056 9908 10090 9942
rect 10128 9908 10162 9942
rect 10200 9908 10234 9942
rect 10272 9908 10306 9942
rect 10344 9908 10378 9942
rect 10416 9908 10450 9942
rect 10488 9908 10522 9942
rect 10560 9908 10594 9942
rect 10632 9908 10666 9942
rect 10704 9908 10738 9942
rect 10776 9908 10810 9942
rect 10848 9908 10882 9942
rect 10920 9908 10954 9942
rect 10992 9908 11026 9942
rect 11064 9908 11098 9942
rect 11136 9908 11170 9942
rect 11208 9908 11242 9942
rect 11280 9908 11314 9942
rect 11352 9908 11386 9942
rect 11424 9908 11458 9942
rect 11496 9908 11530 9942
rect 11568 9908 11602 9942
rect 11640 9908 11674 9942
rect 11712 9908 11746 9942
rect 11784 9908 11818 9942
rect 11856 9908 11890 9942
rect 11928 9908 11962 9942
rect 12000 9908 12034 9942
rect 12072 9908 12106 9942
rect 12144 9908 12178 9942
rect 12216 9908 12250 9942
rect 12288 9908 12322 9942
rect 12360 9908 12394 9942
rect 12432 9908 12466 9942
rect 12504 9908 12538 9942
rect 12576 9908 12610 9942
rect 12648 9908 12682 9942
rect 12720 9908 12754 9942
rect 12792 9908 12826 9942
rect 12864 9908 12898 9942
rect 12936 9908 12970 9942
rect 13008 9908 13042 9942
rect 13080 9908 13114 9942
rect 13152 9908 13186 9942
rect 13224 9908 13258 9942
rect 13296 9908 13330 9942
rect 13368 9908 13402 9942
rect 13440 9908 13474 9942
rect 13512 9908 13546 9942
rect 13584 9908 13618 9942
rect 13656 9908 13690 9942
rect 13728 9908 13762 9942
rect 13800 9908 13834 9942
rect 13872 9908 13906 9942
rect 13944 9908 13978 9942
rect 14016 9908 14050 9942
rect 883 9741 909 9774
rect 909 9741 917 9774
rect 955 9741 977 9774
rect 977 9741 989 9774
rect 1027 9741 1045 9774
rect 1045 9741 1061 9774
rect 1099 9741 1113 9774
rect 1113 9741 1133 9774
rect 1171 9741 1181 9774
rect 1181 9741 1205 9774
rect 1243 9741 1249 9774
rect 1249 9741 1277 9774
rect 1315 9741 1317 9774
rect 1317 9741 1349 9774
rect 1387 9741 1419 9774
rect 1419 9741 1421 9774
rect 1459 9741 1487 9774
rect 1487 9741 1493 9774
rect 1531 9741 1555 9774
rect 1555 9741 1565 9774
rect 1603 9741 1623 9774
rect 1623 9741 1637 9774
rect 1675 9741 1691 9774
rect 1691 9741 1709 9774
rect 1747 9741 1759 9774
rect 1759 9741 1781 9774
rect 1819 9741 1827 9774
rect 1827 9741 1853 9774
rect 1891 9741 1895 9774
rect 1895 9741 1925 9774
rect 883 9740 917 9741
rect 955 9740 989 9741
rect 1027 9740 1061 9741
rect 1099 9740 1133 9741
rect 1171 9740 1205 9741
rect 1243 9740 1277 9741
rect 1315 9740 1349 9741
rect 1387 9740 1421 9741
rect 1459 9740 1493 9741
rect 1531 9740 1565 9741
rect 1603 9740 1637 9741
rect 1675 9740 1709 9741
rect 1747 9740 1781 9741
rect 1819 9740 1853 9741
rect 1891 9740 1925 9741
rect 1963 9740 1997 9774
rect 2035 9741 2065 9774
rect 2065 9741 2069 9774
rect 12883 9741 12911 9774
rect 12911 9741 12917 9774
rect 12955 9741 12979 9774
rect 12979 9741 12989 9774
rect 13027 9741 13047 9774
rect 13047 9741 13061 9774
rect 13099 9741 13115 9774
rect 13115 9741 13133 9774
rect 13171 9741 13183 9774
rect 13183 9741 13205 9774
rect 13243 9741 13251 9774
rect 13251 9741 13277 9774
rect 13315 9741 13319 9774
rect 13319 9741 13349 9774
rect 2035 9740 2069 9741
rect 12883 9740 12917 9741
rect 12955 9740 12989 9741
rect 13027 9740 13061 9741
rect 13099 9740 13133 9741
rect 13171 9740 13205 9741
rect 13243 9740 13277 9741
rect 13315 9740 13349 9741
rect 13387 9740 13421 9774
rect 13459 9741 13489 9774
rect 13489 9741 13493 9774
rect 13531 9741 13557 9774
rect 13557 9741 13565 9774
rect 13603 9741 13625 9774
rect 13625 9741 13637 9774
rect 13675 9741 13693 9774
rect 13693 9741 13709 9774
rect 13747 9741 13761 9774
rect 13761 9741 13781 9774
rect 13819 9741 13829 9774
rect 13829 9741 13853 9774
rect 13891 9741 13897 9774
rect 13897 9741 13925 9774
rect 13963 9741 13965 9774
rect 13965 9741 13997 9774
rect 14035 9741 14067 9774
rect 14067 9741 14069 9774
rect 13459 9740 13493 9741
rect 13531 9740 13565 9741
rect 13603 9740 13637 9741
rect 13675 9740 13709 9741
rect 13747 9740 13781 9741
rect 13819 9740 13853 9741
rect 13891 9740 13925 9741
rect 13963 9740 13997 9741
rect 14035 9740 14069 9741
rect 14614 36157 14643 36190
rect 14643 36157 14648 36190
rect 14614 36156 14648 36157
rect 14614 36089 14643 36118
rect 14643 36089 14648 36118
rect 14614 36084 14648 36089
rect 14614 36021 14643 36046
rect 14643 36021 14648 36046
rect 14614 36012 14648 36021
rect 14614 35953 14643 35974
rect 14643 35953 14648 35974
rect 14614 35940 14648 35953
rect 14614 35885 14643 35902
rect 14643 35885 14648 35902
rect 14614 35868 14648 35885
rect 14614 35817 14643 35830
rect 14643 35817 14648 35830
rect 14614 35796 14648 35817
rect 14614 35749 14643 35758
rect 14643 35749 14648 35758
rect 14614 35724 14648 35749
rect 14614 35681 14643 35686
rect 14643 35681 14648 35686
rect 14614 35652 14648 35681
rect 14614 35613 14643 35614
rect 14643 35613 14648 35614
rect 14614 35580 14648 35613
rect 14614 35511 14648 35542
rect 14614 35508 14643 35511
rect 14643 35508 14648 35511
rect 14614 35443 14648 35470
rect 14614 35436 14643 35443
rect 14643 35436 14648 35443
rect 14614 35375 14648 35398
rect 14614 35364 14643 35375
rect 14643 35364 14648 35375
rect 14614 35307 14648 35326
rect 14614 35292 14643 35307
rect 14643 35292 14648 35307
rect 14614 35239 14648 35254
rect 14614 35220 14643 35239
rect 14643 35220 14648 35239
rect 14614 35171 14648 35182
rect 14614 35148 14643 35171
rect 14643 35148 14648 35171
rect 14614 35103 14648 35110
rect 14614 35076 14643 35103
rect 14643 35076 14648 35103
rect 14614 35035 14648 35038
rect 14614 35004 14643 35035
rect 14643 35004 14648 35035
rect 14614 34933 14643 34966
rect 14643 34933 14648 34966
rect 14614 34932 14648 34933
rect 14614 34865 14643 34894
rect 14643 34865 14648 34894
rect 14614 34860 14648 34865
rect 14614 34797 14643 34822
rect 14643 34797 14648 34822
rect 14614 34788 14648 34797
rect 14614 34729 14643 34750
rect 14643 34729 14648 34750
rect 14614 34716 14648 34729
rect 14614 34661 14643 34678
rect 14643 34661 14648 34678
rect 14614 34644 14648 34661
rect 14614 34593 14643 34606
rect 14643 34593 14648 34606
rect 14614 34572 14648 34593
rect 14614 34525 14643 34534
rect 14643 34525 14648 34534
rect 14614 34500 14648 34525
rect 14614 34457 14643 34462
rect 14643 34457 14648 34462
rect 14614 34428 14648 34457
rect 14614 34389 14643 34390
rect 14643 34389 14648 34390
rect 14614 34356 14648 34389
rect 14614 34287 14648 34318
rect 14614 34284 14643 34287
rect 14643 34284 14648 34287
rect 14614 34219 14648 34246
rect 14614 34212 14643 34219
rect 14643 34212 14648 34219
rect 14614 34151 14648 34174
rect 14614 34140 14643 34151
rect 14643 34140 14648 34151
rect 14614 34083 14648 34102
rect 14614 34068 14643 34083
rect 14643 34068 14648 34083
rect 14614 34015 14648 34030
rect 14614 33996 14643 34015
rect 14643 33996 14648 34015
rect 14614 33947 14648 33958
rect 14614 33924 14643 33947
rect 14643 33924 14648 33947
rect 14614 33879 14648 33886
rect 14614 33852 14643 33879
rect 14643 33852 14648 33879
rect 14614 33811 14648 33814
rect 14614 33780 14643 33811
rect 14643 33780 14648 33811
rect 14614 33709 14643 33742
rect 14643 33709 14648 33742
rect 14614 33708 14648 33709
rect 14614 33641 14643 33670
rect 14643 33641 14648 33670
rect 14614 33636 14648 33641
rect 14614 33573 14643 33598
rect 14643 33573 14648 33598
rect 14614 33564 14648 33573
rect 14614 33505 14643 33526
rect 14643 33505 14648 33526
rect 14614 33492 14648 33505
rect 14614 33437 14643 33454
rect 14643 33437 14648 33454
rect 14614 33420 14648 33437
rect 14614 33369 14643 33382
rect 14643 33369 14648 33382
rect 14614 33348 14648 33369
rect 14614 33301 14643 33310
rect 14643 33301 14648 33310
rect 14614 33276 14648 33301
rect 14614 33233 14643 33238
rect 14643 33233 14648 33238
rect 14614 33204 14648 33233
rect 14614 33165 14643 33166
rect 14643 33165 14648 33166
rect 14614 33132 14648 33165
rect 14614 33063 14648 33094
rect 14614 33060 14643 33063
rect 14643 33060 14648 33063
rect 14614 32995 14648 33022
rect 14614 32988 14643 32995
rect 14643 32988 14648 32995
rect 14614 32927 14648 32950
rect 14614 32916 14643 32927
rect 14643 32916 14648 32927
rect 14614 32859 14648 32878
rect 14614 32844 14643 32859
rect 14643 32844 14648 32859
rect 14614 32791 14648 32806
rect 14614 32772 14643 32791
rect 14643 32772 14648 32791
rect 14614 32723 14648 32734
rect 14614 32700 14643 32723
rect 14643 32700 14648 32723
rect 14614 32655 14648 32662
rect 14614 32628 14643 32655
rect 14643 32628 14648 32655
rect 14614 32587 14648 32590
rect 14614 32556 14643 32587
rect 14643 32556 14648 32587
rect 14614 32485 14643 32518
rect 14643 32485 14648 32518
rect 14614 32484 14648 32485
rect 14614 32417 14643 32446
rect 14643 32417 14648 32446
rect 14614 32412 14648 32417
rect 14614 32349 14643 32374
rect 14643 32349 14648 32374
rect 14614 32340 14648 32349
rect 14614 32281 14643 32302
rect 14643 32281 14648 32302
rect 14614 32268 14648 32281
rect 14614 32213 14643 32230
rect 14643 32213 14648 32230
rect 14614 32196 14648 32213
rect 14614 32145 14643 32158
rect 14643 32145 14648 32158
rect 14614 32124 14648 32145
rect 14614 32077 14643 32086
rect 14643 32077 14648 32086
rect 14614 32052 14648 32077
rect 14614 32009 14643 32014
rect 14643 32009 14648 32014
rect 14614 31980 14648 32009
rect 14614 31941 14643 31942
rect 14643 31941 14648 31942
rect 14614 31908 14648 31941
rect 14614 31839 14648 31870
rect 14614 31836 14643 31839
rect 14643 31836 14648 31839
rect 14614 31771 14648 31798
rect 14614 31764 14643 31771
rect 14643 31764 14648 31771
rect 14614 31703 14648 31726
rect 14614 31692 14643 31703
rect 14643 31692 14648 31703
rect 14614 31635 14648 31654
rect 14614 31620 14643 31635
rect 14643 31620 14648 31635
rect 14614 31567 14648 31582
rect 14614 31548 14643 31567
rect 14643 31548 14648 31567
rect 14614 31499 14648 31510
rect 14614 31476 14643 31499
rect 14643 31476 14648 31499
rect 14614 31431 14648 31438
rect 14614 31404 14643 31431
rect 14643 31404 14648 31431
rect 14614 31363 14648 31366
rect 14614 31332 14643 31363
rect 14643 31332 14648 31363
rect 14614 31261 14643 31294
rect 14643 31261 14648 31294
rect 14614 31260 14648 31261
rect 14614 31193 14643 31222
rect 14643 31193 14648 31222
rect 14614 31188 14648 31193
rect 14614 31125 14643 31150
rect 14643 31125 14648 31150
rect 14614 31116 14648 31125
rect 14614 31057 14643 31078
rect 14643 31057 14648 31078
rect 14614 31044 14648 31057
rect 14614 30989 14643 31006
rect 14643 30989 14648 31006
rect 14614 30972 14648 30989
rect 14614 30921 14643 30934
rect 14643 30921 14648 30934
rect 14614 30900 14648 30921
rect 14614 30853 14643 30862
rect 14643 30853 14648 30862
rect 14614 30828 14648 30853
rect 14614 30785 14643 30790
rect 14643 30785 14648 30790
rect 14614 30756 14648 30785
rect 14614 30717 14643 30718
rect 14643 30717 14648 30718
rect 14614 30684 14648 30717
rect 14614 30615 14648 30646
rect 14614 30612 14643 30615
rect 14643 30612 14648 30615
rect 14614 30547 14648 30574
rect 14614 30540 14643 30547
rect 14643 30540 14648 30547
rect 14614 30479 14648 30502
rect 14614 30468 14643 30479
rect 14643 30468 14648 30479
rect 14614 30411 14648 30430
rect 14614 30396 14643 30411
rect 14643 30396 14648 30411
rect 14614 30343 14648 30358
rect 14614 30324 14643 30343
rect 14643 30324 14648 30343
rect 14614 30275 14648 30286
rect 14614 30252 14643 30275
rect 14643 30252 14648 30275
rect 14614 30207 14648 30214
rect 14614 30180 14643 30207
rect 14643 30180 14648 30207
rect 14614 30139 14648 30142
rect 14614 30108 14643 30139
rect 14643 30108 14648 30139
rect 14614 30037 14643 30070
rect 14643 30037 14648 30070
rect 14614 30036 14648 30037
rect 14614 29969 14643 29998
rect 14643 29969 14648 29998
rect 14614 29964 14648 29969
rect 14614 29901 14643 29926
rect 14643 29901 14648 29926
rect 14614 29892 14648 29901
rect 14614 29833 14643 29854
rect 14643 29833 14648 29854
rect 14614 29820 14648 29833
rect 14614 29765 14643 29782
rect 14643 29765 14648 29782
rect 14614 29748 14648 29765
rect 14614 29697 14643 29710
rect 14643 29697 14648 29710
rect 14614 29676 14648 29697
rect 14614 29629 14643 29638
rect 14643 29629 14648 29638
rect 14614 29604 14648 29629
rect 14614 29561 14643 29566
rect 14643 29561 14648 29566
rect 14614 29532 14648 29561
rect 14614 29493 14643 29494
rect 14643 29493 14648 29494
rect 14614 29460 14648 29493
rect 14614 29391 14648 29422
rect 14614 29388 14643 29391
rect 14643 29388 14648 29391
rect 14614 29323 14648 29350
rect 14614 29316 14643 29323
rect 14643 29316 14648 29323
rect 14614 29255 14648 29278
rect 14614 29244 14643 29255
rect 14643 29244 14648 29255
rect 14614 29187 14648 29206
rect 14614 29172 14643 29187
rect 14643 29172 14648 29187
rect 14614 29119 14648 29134
rect 14614 29100 14643 29119
rect 14643 29100 14648 29119
rect 14614 29051 14648 29062
rect 14614 29028 14643 29051
rect 14643 29028 14648 29051
rect 14614 28983 14648 28990
rect 14614 28956 14643 28983
rect 14643 28956 14648 28983
rect 14614 28915 14648 28918
rect 14614 28884 14643 28915
rect 14643 28884 14648 28915
rect 14614 28813 14643 28846
rect 14643 28813 14648 28846
rect 14614 28812 14648 28813
rect 14614 28745 14643 28774
rect 14643 28745 14648 28774
rect 14614 28740 14648 28745
rect 14614 28677 14643 28702
rect 14643 28677 14648 28702
rect 14614 28668 14648 28677
rect 14614 28609 14643 28630
rect 14643 28609 14648 28630
rect 14614 28596 14648 28609
rect 14614 28541 14643 28558
rect 14643 28541 14648 28558
rect 14614 28524 14648 28541
rect 14614 28473 14643 28486
rect 14643 28473 14648 28486
rect 14614 28452 14648 28473
rect 14614 28405 14643 28414
rect 14643 28405 14648 28414
rect 14614 28380 14648 28405
rect 14614 28337 14643 28342
rect 14643 28337 14648 28342
rect 14614 28308 14648 28337
rect 14614 28269 14643 28270
rect 14643 28269 14648 28270
rect 14614 28236 14648 28269
rect 14614 28167 14648 28198
rect 14614 28164 14643 28167
rect 14643 28164 14648 28167
rect 14614 28099 14648 28126
rect 14614 28092 14643 28099
rect 14643 28092 14648 28099
rect 14614 28031 14648 28054
rect 14614 28020 14643 28031
rect 14643 28020 14648 28031
rect 14614 27963 14648 27982
rect 14614 27948 14643 27963
rect 14643 27948 14648 27963
rect 14614 27895 14648 27910
rect 14614 27876 14643 27895
rect 14643 27876 14648 27895
rect 14614 27827 14648 27838
rect 14614 27804 14643 27827
rect 14643 27804 14648 27827
rect 14614 27759 14648 27766
rect 14614 27732 14643 27759
rect 14643 27732 14648 27759
rect 14614 27691 14648 27694
rect 14614 27660 14643 27691
rect 14643 27660 14648 27691
rect 14614 27589 14643 27622
rect 14643 27589 14648 27622
rect 14614 27588 14648 27589
rect 14614 27521 14643 27550
rect 14643 27521 14648 27550
rect 14614 27516 14648 27521
rect 14614 27453 14643 27478
rect 14643 27453 14648 27478
rect 14614 27444 14648 27453
rect 14614 27385 14643 27406
rect 14643 27385 14648 27406
rect 14614 27372 14648 27385
rect 14614 27317 14643 27334
rect 14643 27317 14648 27334
rect 14614 27300 14648 27317
rect 14614 27249 14643 27262
rect 14643 27249 14648 27262
rect 14614 27228 14648 27249
rect 14614 27181 14643 27190
rect 14643 27181 14648 27190
rect 14614 27156 14648 27181
rect 14614 27113 14643 27118
rect 14643 27113 14648 27118
rect 14614 27084 14648 27113
rect 14614 27045 14643 27046
rect 14643 27045 14648 27046
rect 14614 27012 14648 27045
rect 14614 26943 14648 26974
rect 14614 26940 14643 26943
rect 14643 26940 14648 26943
rect 14614 26875 14648 26902
rect 14614 26868 14643 26875
rect 14643 26868 14648 26875
rect 14614 26807 14648 26830
rect 14614 26796 14643 26807
rect 14643 26796 14648 26807
rect 14614 26739 14648 26758
rect 14614 26724 14643 26739
rect 14643 26724 14648 26739
rect 14614 26671 14648 26686
rect 14614 26652 14643 26671
rect 14643 26652 14648 26671
rect 14614 26603 14648 26614
rect 14614 26580 14643 26603
rect 14643 26580 14648 26603
rect 14614 26535 14648 26542
rect 14614 26508 14643 26535
rect 14643 26508 14648 26535
rect 14614 26467 14648 26470
rect 14614 26436 14643 26467
rect 14643 26436 14648 26467
rect 14614 26365 14643 26398
rect 14643 26365 14648 26398
rect 14614 26364 14648 26365
rect 14614 26297 14643 26326
rect 14643 26297 14648 26326
rect 14614 26292 14648 26297
rect 14614 26229 14643 26254
rect 14643 26229 14648 26254
rect 14614 26220 14648 26229
rect 14614 26161 14643 26182
rect 14643 26161 14648 26182
rect 14614 26148 14648 26161
rect 14614 26093 14643 26110
rect 14643 26093 14648 26110
rect 14614 26076 14648 26093
rect 14614 26025 14643 26038
rect 14643 26025 14648 26038
rect 14614 26004 14648 26025
rect 14614 25957 14643 25966
rect 14643 25957 14648 25966
rect 14614 25932 14648 25957
rect 14614 25889 14643 25894
rect 14643 25889 14648 25894
rect 14614 25860 14648 25889
rect 14614 25821 14643 25822
rect 14643 25821 14648 25822
rect 14614 25788 14648 25821
rect 14614 25719 14648 25750
rect 14614 25716 14643 25719
rect 14643 25716 14648 25719
rect 14614 25651 14648 25678
rect 14614 25644 14643 25651
rect 14643 25644 14648 25651
rect 14614 25583 14648 25606
rect 14614 25572 14643 25583
rect 14643 25572 14648 25583
rect 14614 25515 14648 25534
rect 14614 25500 14643 25515
rect 14643 25500 14648 25515
rect 14614 25447 14648 25462
rect 14614 25428 14643 25447
rect 14643 25428 14648 25447
rect 14614 25379 14648 25390
rect 14614 25356 14643 25379
rect 14643 25356 14648 25379
rect 14614 25311 14648 25318
rect 14614 25284 14643 25311
rect 14643 25284 14648 25311
rect 14614 25243 14648 25246
rect 14614 25212 14643 25243
rect 14643 25212 14648 25243
rect 14614 25141 14643 25174
rect 14643 25141 14648 25174
rect 14614 25140 14648 25141
rect 14614 25073 14643 25102
rect 14643 25073 14648 25102
rect 14614 25068 14648 25073
rect 14614 25005 14643 25030
rect 14643 25005 14648 25030
rect 14614 24996 14648 25005
rect 14614 24937 14643 24958
rect 14643 24937 14648 24958
rect 14614 24924 14648 24937
rect 14614 24869 14643 24886
rect 14643 24869 14648 24886
rect 14614 24852 14648 24869
rect 14614 24801 14643 24814
rect 14643 24801 14648 24814
rect 14614 24780 14648 24801
rect 14614 24733 14643 24742
rect 14643 24733 14648 24742
rect 14614 24708 14648 24733
rect 14614 24665 14643 24670
rect 14643 24665 14648 24670
rect 14614 24636 14648 24665
rect 14614 24597 14643 24598
rect 14643 24597 14648 24598
rect 14614 24564 14648 24597
rect 14614 24495 14648 24526
rect 14614 24492 14643 24495
rect 14643 24492 14648 24495
rect 14614 24427 14648 24454
rect 14614 24420 14643 24427
rect 14643 24420 14648 24427
rect 14614 24359 14648 24382
rect 14614 24348 14643 24359
rect 14643 24348 14648 24359
rect 14614 24291 14648 24310
rect 14614 24276 14643 24291
rect 14643 24276 14648 24291
rect 14614 24223 14648 24238
rect 14614 24204 14643 24223
rect 14643 24204 14648 24223
rect 14614 24155 14648 24166
rect 14614 24132 14643 24155
rect 14643 24132 14648 24155
rect 14614 24087 14648 24094
rect 14614 24060 14643 24087
rect 14643 24060 14648 24087
rect 14614 24019 14648 24022
rect 14614 23988 14643 24019
rect 14643 23988 14648 24019
rect 14614 23917 14643 23950
rect 14643 23917 14648 23950
rect 14614 23916 14648 23917
rect 14614 23849 14643 23878
rect 14643 23849 14648 23878
rect 14614 23844 14648 23849
rect 14614 23781 14643 23806
rect 14643 23781 14648 23806
rect 14614 23772 14648 23781
rect 14614 23713 14643 23734
rect 14643 23713 14648 23734
rect 14614 23700 14648 23713
rect 14614 23645 14643 23662
rect 14643 23645 14648 23662
rect 14614 23628 14648 23645
rect 14614 23577 14643 23590
rect 14643 23577 14648 23590
rect 14614 23556 14648 23577
rect 14614 23509 14643 23518
rect 14643 23509 14648 23518
rect 14614 23484 14648 23509
rect 14614 23441 14643 23446
rect 14643 23441 14648 23446
rect 14614 23412 14648 23441
rect 14614 23373 14643 23374
rect 14643 23373 14648 23374
rect 14614 23340 14648 23373
rect 14614 23271 14648 23302
rect 14614 23268 14643 23271
rect 14643 23268 14648 23271
rect 14614 23203 14648 23230
rect 14614 23196 14643 23203
rect 14643 23196 14648 23203
rect 14614 23135 14648 23158
rect 14614 23124 14643 23135
rect 14643 23124 14648 23135
rect 14614 23067 14648 23086
rect 14614 23052 14643 23067
rect 14643 23052 14648 23067
rect 14614 22999 14648 23014
rect 14614 22980 14643 22999
rect 14643 22980 14648 22999
rect 14614 22931 14648 22942
rect 14614 22908 14643 22931
rect 14643 22908 14648 22931
rect 14614 22863 14648 22870
rect 14614 22836 14643 22863
rect 14643 22836 14648 22863
rect 14614 22795 14648 22798
rect 14614 22764 14643 22795
rect 14643 22764 14648 22795
rect 14614 22693 14643 22726
rect 14643 22693 14648 22726
rect 14614 22692 14648 22693
rect 14614 22625 14643 22654
rect 14643 22625 14648 22654
rect 14614 22620 14648 22625
rect 14614 22557 14643 22582
rect 14643 22557 14648 22582
rect 14614 22548 14648 22557
rect 14614 22489 14643 22510
rect 14643 22489 14648 22510
rect 14614 22476 14648 22489
rect 14614 22421 14643 22438
rect 14643 22421 14648 22438
rect 14614 22404 14648 22421
rect 14614 22353 14643 22366
rect 14643 22353 14648 22366
rect 14614 22332 14648 22353
rect 14614 22285 14643 22294
rect 14643 22285 14648 22294
rect 14614 22260 14648 22285
rect 14614 22217 14643 22222
rect 14643 22217 14648 22222
rect 14614 22188 14648 22217
rect 14614 22149 14643 22150
rect 14643 22149 14648 22150
rect 14614 22116 14648 22149
rect 14614 22047 14648 22078
rect 14614 22044 14643 22047
rect 14643 22044 14648 22047
rect 14614 21979 14648 22006
rect 14614 21972 14643 21979
rect 14643 21972 14648 21979
rect 14614 21911 14648 21934
rect 14614 21900 14643 21911
rect 14643 21900 14648 21911
rect 14614 21843 14648 21862
rect 14614 21828 14643 21843
rect 14643 21828 14648 21843
rect 14614 21775 14648 21790
rect 14614 21756 14643 21775
rect 14643 21756 14648 21775
rect 14614 21707 14648 21718
rect 14614 21684 14643 21707
rect 14643 21684 14648 21707
rect 14614 21639 14648 21646
rect 14614 21612 14643 21639
rect 14643 21612 14648 21639
rect 14614 21571 14648 21574
rect 14614 21540 14643 21571
rect 14643 21540 14648 21571
rect 14614 21469 14643 21502
rect 14643 21469 14648 21502
rect 14614 21468 14648 21469
rect 14614 21401 14643 21430
rect 14643 21401 14648 21430
rect 14614 21396 14648 21401
rect 14614 21333 14643 21358
rect 14643 21333 14648 21358
rect 14614 21324 14648 21333
rect 14614 21265 14643 21286
rect 14643 21265 14648 21286
rect 14614 21252 14648 21265
rect 14614 21197 14643 21214
rect 14643 21197 14648 21214
rect 14614 21180 14648 21197
rect 14614 21129 14643 21142
rect 14643 21129 14648 21142
rect 14614 21108 14648 21129
rect 14614 21061 14643 21070
rect 14643 21061 14648 21070
rect 14614 21036 14648 21061
rect 14614 20993 14643 20998
rect 14643 20993 14648 20998
rect 14614 20964 14648 20993
rect 14614 20925 14643 20926
rect 14643 20925 14648 20926
rect 14614 20892 14648 20925
rect 14614 20823 14648 20854
rect 14614 20820 14643 20823
rect 14643 20820 14648 20823
rect 14614 20755 14648 20782
rect 14614 20748 14643 20755
rect 14643 20748 14648 20755
rect 14614 20687 14648 20710
rect 14614 20676 14643 20687
rect 14643 20676 14648 20687
rect 14614 20619 14648 20638
rect 14614 20604 14643 20619
rect 14643 20604 14648 20619
rect 14614 20551 14648 20566
rect 14614 20532 14643 20551
rect 14643 20532 14648 20551
rect 14614 20483 14648 20494
rect 14614 20460 14643 20483
rect 14643 20460 14648 20483
rect 14614 20415 14648 20422
rect 14614 20388 14643 20415
rect 14643 20388 14648 20415
rect 14614 20347 14648 20350
rect 14614 20316 14643 20347
rect 14643 20316 14648 20347
rect 14614 20245 14643 20278
rect 14643 20245 14648 20278
rect 14614 20244 14648 20245
rect 14614 20177 14643 20206
rect 14643 20177 14648 20206
rect 14614 20172 14648 20177
rect 14614 20109 14643 20134
rect 14643 20109 14648 20134
rect 14614 20100 14648 20109
rect 14614 20041 14643 20062
rect 14643 20041 14648 20062
rect 14614 20028 14648 20041
rect 14614 19973 14643 19990
rect 14643 19973 14648 19990
rect 14614 19956 14648 19973
rect 14614 19905 14643 19918
rect 14643 19905 14648 19918
rect 14614 19884 14648 19905
rect 14614 19837 14643 19846
rect 14643 19837 14648 19846
rect 14614 19812 14648 19837
rect 14614 19769 14643 19774
rect 14643 19769 14648 19774
rect 14614 19740 14648 19769
rect 14614 19701 14643 19702
rect 14643 19701 14648 19702
rect 14614 19668 14648 19701
rect 14614 19599 14648 19630
rect 14614 19596 14643 19599
rect 14643 19596 14648 19599
rect 14614 19531 14648 19558
rect 14614 19524 14643 19531
rect 14643 19524 14648 19531
rect 14614 19463 14648 19486
rect 14614 19452 14643 19463
rect 14643 19452 14648 19463
rect 14614 19395 14648 19414
rect 14614 19380 14643 19395
rect 14643 19380 14648 19395
rect 14614 19327 14648 19342
rect 14614 19308 14643 19327
rect 14643 19308 14648 19327
rect 14614 19259 14648 19270
rect 14614 19236 14643 19259
rect 14643 19236 14648 19259
rect 14614 19191 14648 19198
rect 14614 19164 14643 19191
rect 14643 19164 14648 19191
rect 14614 19123 14648 19126
rect 14614 19092 14643 19123
rect 14643 19092 14648 19123
rect 14614 19021 14643 19054
rect 14643 19021 14648 19054
rect 14614 19020 14648 19021
rect 14614 18953 14643 18982
rect 14643 18953 14648 18982
rect 14614 18948 14648 18953
rect 14614 18885 14643 18910
rect 14643 18885 14648 18910
rect 14614 18876 14648 18885
rect 14614 18817 14643 18838
rect 14643 18817 14648 18838
rect 14614 18804 14648 18817
rect 14614 18749 14643 18766
rect 14643 18749 14648 18766
rect 14614 18732 14648 18749
rect 14614 18681 14643 18694
rect 14643 18681 14648 18694
rect 14614 18660 14648 18681
rect 14614 18613 14643 18622
rect 14643 18613 14648 18622
rect 14614 18588 14648 18613
rect 14614 18545 14643 18550
rect 14643 18545 14648 18550
rect 14614 18516 14648 18545
rect 14614 18477 14643 18478
rect 14643 18477 14648 18478
rect 14614 18444 14648 18477
rect 14614 18375 14648 18406
rect 14614 18372 14643 18375
rect 14643 18372 14648 18375
rect 14614 18307 14648 18334
rect 14614 18300 14643 18307
rect 14643 18300 14648 18307
rect 14614 18239 14648 18262
rect 14614 18228 14643 18239
rect 14643 18228 14648 18239
rect 14614 18171 14648 18190
rect 14614 18156 14643 18171
rect 14643 18156 14648 18171
rect 14614 18103 14648 18118
rect 14614 18084 14643 18103
rect 14643 18084 14648 18103
rect 14614 18035 14648 18046
rect 14614 18012 14643 18035
rect 14643 18012 14648 18035
rect 14614 17967 14648 17974
rect 14614 17940 14643 17967
rect 14643 17940 14648 17967
rect 14614 17899 14648 17902
rect 14614 17868 14643 17899
rect 14643 17868 14648 17899
rect 14614 17797 14643 17830
rect 14643 17797 14648 17830
rect 14614 17796 14648 17797
rect 14614 17729 14643 17758
rect 14643 17729 14648 17758
rect 14614 17724 14648 17729
rect 14614 17661 14643 17686
rect 14643 17661 14648 17686
rect 14614 17652 14648 17661
rect 14614 17593 14643 17614
rect 14643 17593 14648 17614
rect 14614 17580 14648 17593
rect 14614 17525 14643 17542
rect 14643 17525 14648 17542
rect 14614 17508 14648 17525
rect 14614 17457 14643 17470
rect 14643 17457 14648 17470
rect 14614 17436 14648 17457
rect 14614 17389 14643 17398
rect 14643 17389 14648 17398
rect 14614 17364 14648 17389
rect 14614 17321 14643 17326
rect 14643 17321 14648 17326
rect 14614 17292 14648 17321
rect 14614 17253 14643 17254
rect 14643 17253 14648 17254
rect 14614 17220 14648 17253
rect 14614 17151 14648 17182
rect 14614 17148 14643 17151
rect 14643 17148 14648 17151
rect 14614 17083 14648 17110
rect 14614 17076 14643 17083
rect 14643 17076 14648 17083
rect 14614 17015 14648 17038
rect 14614 17004 14643 17015
rect 14643 17004 14648 17015
rect 14614 16947 14648 16966
rect 14614 16932 14643 16947
rect 14643 16932 14648 16947
rect 14614 16879 14648 16894
rect 14614 16860 14643 16879
rect 14643 16860 14648 16879
rect 14614 16811 14648 16822
rect 14614 16788 14643 16811
rect 14643 16788 14648 16811
rect 14614 16743 14648 16750
rect 14614 16716 14643 16743
rect 14643 16716 14648 16743
rect 14614 16675 14648 16678
rect 14614 16644 14643 16675
rect 14643 16644 14648 16675
rect 14614 16573 14643 16606
rect 14643 16573 14648 16606
rect 14614 16572 14648 16573
rect 14614 16505 14643 16534
rect 14643 16505 14648 16534
rect 14614 16500 14648 16505
rect 14614 16437 14643 16462
rect 14643 16437 14648 16462
rect 14614 16428 14648 16437
rect 14614 16369 14643 16390
rect 14643 16369 14648 16390
rect 14614 16356 14648 16369
rect 14614 16301 14643 16318
rect 14643 16301 14648 16318
rect 14614 16284 14648 16301
rect 14614 16233 14643 16246
rect 14643 16233 14648 16246
rect 14614 16212 14648 16233
rect 14614 16165 14643 16174
rect 14643 16165 14648 16174
rect 14614 16140 14648 16165
rect 14614 16097 14643 16102
rect 14643 16097 14648 16102
rect 14614 16068 14648 16097
rect 14614 16029 14643 16030
rect 14643 16029 14648 16030
rect 14614 15996 14648 16029
rect 14614 15927 14648 15958
rect 14614 15924 14643 15927
rect 14643 15924 14648 15927
rect 14614 15859 14648 15886
rect 14614 15852 14643 15859
rect 14643 15852 14648 15859
rect 14614 15791 14648 15814
rect 14614 15780 14643 15791
rect 14643 15780 14648 15791
rect 14614 15723 14648 15742
rect 14614 15708 14643 15723
rect 14643 15708 14648 15723
rect 14614 15655 14648 15670
rect 14614 15636 14643 15655
rect 14643 15636 14648 15655
rect 14614 15587 14648 15598
rect 14614 15564 14643 15587
rect 14643 15564 14648 15587
rect 14614 15519 14648 15526
rect 14614 15492 14643 15519
rect 14643 15492 14648 15519
rect 14614 15451 14648 15454
rect 14614 15420 14643 15451
rect 14643 15420 14648 15451
rect 14614 15349 14643 15382
rect 14643 15349 14648 15382
rect 14614 15348 14648 15349
rect 14614 15281 14643 15310
rect 14643 15281 14648 15310
rect 14614 15276 14648 15281
rect 14614 15213 14643 15238
rect 14643 15213 14648 15238
rect 14614 15204 14648 15213
rect 14614 15145 14643 15166
rect 14643 15145 14648 15166
rect 14614 15132 14648 15145
rect 14614 15077 14643 15094
rect 14643 15077 14648 15094
rect 14614 15060 14648 15077
rect 14614 15009 14643 15022
rect 14643 15009 14648 15022
rect 14614 14988 14648 15009
rect 14614 14941 14643 14950
rect 14643 14941 14648 14950
rect 14614 14916 14648 14941
rect 14614 14873 14643 14878
rect 14643 14873 14648 14878
rect 14614 14844 14648 14873
rect 14614 14805 14643 14806
rect 14643 14805 14648 14806
rect 14614 14772 14648 14805
rect 14614 14703 14648 14734
rect 14614 14700 14643 14703
rect 14643 14700 14648 14703
rect 14614 14635 14648 14662
rect 14614 14628 14643 14635
rect 14643 14628 14648 14635
rect 14614 14567 14648 14590
rect 14614 14556 14643 14567
rect 14643 14556 14648 14567
rect 14614 14499 14648 14518
rect 14614 14484 14643 14499
rect 14643 14484 14648 14499
rect 14614 14431 14648 14446
rect 14614 14412 14643 14431
rect 14643 14412 14648 14431
rect 14614 14363 14648 14374
rect 14614 14340 14643 14363
rect 14643 14340 14648 14363
rect 14614 14295 14648 14302
rect 14614 14268 14643 14295
rect 14643 14268 14648 14295
rect 14614 14227 14648 14230
rect 14614 14196 14643 14227
rect 14643 14196 14648 14227
rect 14614 14125 14643 14158
rect 14643 14125 14648 14158
rect 14614 14124 14648 14125
rect 14614 14057 14643 14086
rect 14643 14057 14648 14086
rect 14614 14052 14648 14057
rect 14614 13989 14643 14014
rect 14643 13989 14648 14014
rect 14614 13980 14648 13989
rect 14614 13921 14643 13942
rect 14643 13921 14648 13942
rect 14614 13908 14648 13921
rect 14614 13853 14643 13870
rect 14643 13853 14648 13870
rect 14614 13836 14648 13853
rect 14614 13785 14643 13798
rect 14643 13785 14648 13798
rect 14614 13764 14648 13785
rect 14614 13717 14643 13726
rect 14643 13717 14648 13726
rect 14614 13692 14648 13717
rect 14614 13649 14643 13654
rect 14643 13649 14648 13654
rect 14614 13620 14648 13649
rect 14614 13581 14643 13582
rect 14643 13581 14648 13582
rect 14614 13548 14648 13581
rect 14614 13479 14648 13510
rect 14614 13476 14643 13479
rect 14643 13476 14648 13479
rect 14614 13411 14648 13438
rect 14614 13404 14643 13411
rect 14643 13404 14648 13411
rect 14614 13343 14648 13366
rect 14614 13332 14643 13343
rect 14643 13332 14648 13343
rect 14614 13275 14648 13294
rect 14614 13260 14643 13275
rect 14643 13260 14648 13275
rect 14614 13207 14648 13222
rect 14614 13188 14643 13207
rect 14643 13188 14648 13207
rect 14614 13139 14648 13150
rect 14614 13116 14643 13139
rect 14643 13116 14648 13139
rect 14614 13071 14648 13078
rect 14614 13044 14643 13071
rect 14643 13044 14648 13071
rect 14614 13003 14648 13006
rect 14614 12972 14643 13003
rect 14643 12972 14648 13003
rect 14614 12901 14643 12934
rect 14643 12901 14648 12934
rect 14614 12900 14648 12901
rect 14614 12833 14643 12862
rect 14643 12833 14648 12862
rect 14614 12828 14648 12833
rect 14614 12765 14643 12790
rect 14643 12765 14648 12790
rect 14614 12756 14648 12765
rect 14614 12697 14643 12718
rect 14643 12697 14648 12718
rect 14614 12684 14648 12697
rect 14614 12629 14643 12646
rect 14643 12629 14648 12646
rect 14614 12612 14648 12629
rect 14614 12561 14643 12574
rect 14643 12561 14648 12574
rect 14614 12540 14648 12561
rect 14614 12493 14643 12502
rect 14643 12493 14648 12502
rect 14614 12468 14648 12493
rect 14614 12425 14643 12430
rect 14643 12425 14648 12430
rect 14614 12396 14648 12425
rect 14614 12357 14643 12358
rect 14643 12357 14648 12358
rect 14614 12324 14648 12357
rect 14614 12255 14648 12286
rect 14614 12252 14643 12255
rect 14643 12252 14648 12255
rect 14614 12187 14648 12214
rect 14614 12180 14643 12187
rect 14643 12180 14648 12187
rect 14614 12119 14648 12142
rect 14614 12108 14643 12119
rect 14643 12108 14648 12119
rect 14614 12051 14648 12070
rect 14614 12036 14643 12051
rect 14643 12036 14648 12051
rect 14614 11983 14648 11998
rect 14614 11964 14643 11983
rect 14643 11964 14648 11983
rect 14614 11915 14648 11926
rect 14614 11892 14643 11915
rect 14643 11892 14648 11915
rect 14614 11847 14648 11854
rect 14614 11820 14643 11847
rect 14643 11820 14648 11847
rect 14614 11779 14648 11782
rect 14614 11748 14643 11779
rect 14643 11748 14648 11779
rect 14614 11677 14643 11710
rect 14643 11677 14648 11710
rect 14614 11676 14648 11677
rect 14614 11609 14643 11638
rect 14643 11609 14648 11638
rect 14614 11604 14648 11609
rect 14614 11541 14643 11566
rect 14643 11541 14648 11566
rect 14614 11532 14648 11541
rect 14614 11473 14643 11494
rect 14643 11473 14648 11494
rect 14614 11460 14648 11473
rect 14614 11405 14643 11422
rect 14643 11405 14648 11422
rect 14614 11388 14648 11405
rect 14614 11337 14643 11350
rect 14643 11337 14648 11350
rect 14614 11316 14648 11337
rect 14614 11269 14643 11278
rect 14643 11269 14648 11278
rect 14614 11244 14648 11269
rect 14614 11201 14643 11206
rect 14643 11201 14648 11206
rect 14614 11172 14648 11201
rect 14614 11133 14643 11134
rect 14643 11133 14648 11134
rect 14614 11100 14648 11133
rect 14614 11031 14648 11062
rect 14614 11028 14643 11031
rect 14643 11028 14648 11031
rect 14614 10963 14648 10990
rect 14614 10956 14643 10963
rect 14643 10956 14648 10963
rect 14614 10895 14648 10918
rect 14614 10884 14643 10895
rect 14643 10884 14648 10895
rect 14614 10827 14648 10846
rect 14614 10812 14643 10827
rect 14643 10812 14648 10827
rect 14614 10759 14648 10774
rect 14614 10740 14643 10759
rect 14643 10740 14648 10759
rect 14614 10691 14648 10702
rect 14614 10668 14643 10691
rect 14643 10668 14648 10691
rect 14614 10623 14648 10630
rect 14614 10596 14643 10623
rect 14643 10596 14648 10623
rect 14614 10555 14648 10558
rect 14614 10524 14643 10555
rect 14643 10524 14648 10555
rect 14614 10453 14643 10486
rect 14643 10453 14648 10486
rect 14614 10452 14648 10453
rect 14614 10385 14643 10414
rect 14643 10385 14648 10414
rect 14614 10380 14648 10385
rect 14614 10317 14643 10342
rect 14643 10317 14648 10342
rect 14614 10308 14648 10317
rect 14614 10249 14643 10270
rect 14643 10249 14648 10270
rect 14614 10236 14648 10249
rect 14614 10181 14643 10198
rect 14643 10181 14648 10198
rect 14614 10164 14648 10181
rect 14614 10113 14643 10126
rect 14643 10113 14648 10126
rect 14614 10092 14648 10113
rect 14614 10045 14643 10054
rect 14643 10045 14648 10054
rect 14614 10020 14648 10045
rect 14614 9977 14643 9982
rect 14643 9977 14648 9982
rect 14614 9948 14648 9977
rect 14614 9909 14643 9910
rect 14643 9909 14648 9910
rect 14614 9876 14648 9909
rect 14614 9807 14648 9838
rect 14614 9804 14643 9807
rect 14643 9804 14648 9807
rect 14614 9739 14648 9766
rect 320 9679 354 9697
rect 320 9663 322 9679
rect 322 9663 354 9679
rect 14614 9732 14643 9739
rect 14643 9732 14648 9739
rect 14614 9671 14648 9694
rect 14614 9660 14643 9671
rect 14643 9660 14648 9671
rect 320 9418 354 9452
rect 610 9420 612 9452
rect 612 9420 644 9452
rect 2311 9420 2312 9452
rect 2312 9420 2345 9452
rect 2383 9420 2414 9452
rect 2414 9420 2417 9452
rect 2455 9420 2482 9452
rect 2482 9420 2489 9452
rect 2527 9420 2550 9452
rect 2550 9420 2561 9452
rect 2599 9420 2618 9452
rect 2618 9420 2633 9452
rect 2671 9420 2686 9452
rect 2686 9420 2705 9452
rect 2743 9420 2754 9452
rect 2754 9420 2777 9452
rect 2815 9420 2822 9452
rect 2822 9420 2849 9452
rect 2887 9420 2890 9452
rect 2890 9420 2921 9452
rect 2959 9420 2992 9452
rect 2992 9420 2993 9452
rect 3031 9420 3060 9452
rect 3060 9420 3065 9452
rect 3103 9420 3128 9452
rect 3128 9420 3137 9452
rect 3175 9420 3196 9452
rect 3196 9420 3209 9452
rect 3247 9420 3264 9452
rect 3264 9420 3281 9452
rect 3319 9420 3332 9452
rect 3332 9420 3353 9452
rect 3391 9420 3400 9452
rect 3400 9420 3425 9452
rect 3463 9420 3468 9452
rect 3468 9420 3497 9452
rect 3535 9420 3536 9452
rect 3536 9420 3569 9452
rect 3607 9420 3638 9452
rect 3638 9420 3641 9452
rect 3679 9420 3706 9452
rect 3706 9420 3713 9452
rect 3751 9420 3774 9452
rect 3774 9420 3785 9452
rect 3823 9420 3842 9452
rect 3842 9420 3857 9452
rect 3895 9420 3910 9452
rect 3910 9420 3929 9452
rect 3967 9420 3978 9452
rect 3978 9420 4001 9452
rect 4039 9420 4046 9452
rect 4046 9420 4073 9452
rect 4111 9420 4114 9452
rect 4114 9420 4145 9452
rect 4183 9420 4216 9452
rect 4216 9420 4217 9452
rect 4255 9420 4284 9452
rect 4284 9420 4289 9452
rect 4327 9420 4352 9452
rect 4352 9420 4361 9452
rect 4399 9420 4420 9452
rect 4420 9420 4433 9452
rect 4471 9420 4488 9452
rect 4488 9420 4505 9452
rect 4543 9420 4556 9452
rect 4556 9420 4577 9452
rect 4615 9420 4624 9452
rect 4624 9420 4649 9452
rect 4687 9420 4692 9452
rect 4692 9420 4721 9452
rect 4759 9420 4760 9452
rect 4760 9420 4793 9452
rect 4831 9420 4862 9452
rect 4862 9420 4865 9452
rect 4903 9420 4930 9452
rect 4930 9420 4937 9452
rect 4975 9420 4998 9452
rect 4998 9420 5009 9452
rect 5047 9420 5066 9452
rect 5066 9420 5081 9452
rect 5119 9420 5134 9452
rect 5134 9420 5153 9452
rect 5191 9420 5202 9452
rect 5202 9420 5225 9452
rect 5263 9420 5270 9452
rect 5270 9420 5297 9452
rect 5335 9420 5338 9452
rect 5338 9420 5369 9452
rect 5407 9420 5440 9452
rect 5440 9420 5441 9452
rect 5479 9420 5508 9452
rect 5508 9420 5513 9452
rect 5551 9420 5576 9452
rect 5576 9420 5585 9452
rect 5623 9420 5644 9452
rect 5644 9420 5657 9452
rect 5695 9420 5712 9452
rect 5712 9420 5729 9452
rect 5767 9420 5780 9452
rect 5780 9420 5801 9452
rect 5839 9420 5848 9452
rect 5848 9420 5873 9452
rect 5911 9420 5916 9452
rect 5916 9420 5945 9452
rect 5983 9420 5984 9452
rect 5984 9420 6017 9452
rect 6055 9420 6086 9452
rect 6086 9420 6089 9452
rect 6127 9420 6154 9452
rect 6154 9420 6161 9452
rect 6199 9420 6222 9452
rect 6222 9420 6233 9452
rect 6271 9420 6290 9452
rect 6290 9420 6305 9452
rect 6343 9420 6358 9452
rect 6358 9420 6377 9452
rect 6415 9420 6426 9452
rect 6426 9420 6449 9452
rect 6487 9420 6494 9452
rect 6494 9420 6521 9452
rect 6559 9420 6562 9452
rect 6562 9420 6593 9452
rect 6631 9420 6664 9452
rect 6664 9420 6665 9452
rect 6703 9420 6732 9452
rect 6732 9420 6737 9452
rect 6775 9420 6800 9452
rect 6800 9420 6809 9452
rect 6847 9420 6868 9452
rect 6868 9420 6881 9452
rect 6919 9420 6936 9452
rect 6936 9420 6953 9452
rect 6991 9420 7004 9452
rect 7004 9420 7025 9452
rect 7063 9420 7072 9452
rect 7072 9420 7097 9452
rect 7135 9420 7140 9452
rect 7140 9420 7169 9452
rect 7207 9420 7208 9452
rect 7208 9420 7241 9452
rect 7279 9420 7310 9452
rect 7310 9420 7313 9452
rect 7351 9420 7378 9452
rect 7378 9420 7385 9452
rect 7423 9420 7446 9452
rect 7446 9420 7457 9452
rect 7495 9420 7514 9452
rect 7514 9420 7529 9452
rect 7567 9420 7582 9452
rect 7582 9420 7601 9452
rect 7639 9420 7650 9452
rect 7650 9420 7673 9452
rect 7711 9420 7718 9452
rect 7718 9420 7745 9452
rect 7783 9420 7786 9452
rect 7786 9420 7817 9452
rect 7855 9420 7888 9452
rect 7888 9420 7889 9452
rect 7927 9420 7956 9452
rect 7956 9420 7961 9452
rect 7999 9420 8024 9452
rect 8024 9420 8033 9452
rect 8071 9420 8092 9452
rect 8092 9420 8105 9452
rect 8143 9420 8160 9452
rect 8160 9420 8177 9452
rect 8215 9420 8228 9452
rect 8228 9420 8249 9452
rect 8287 9420 8296 9452
rect 8296 9420 8321 9452
rect 8359 9420 8364 9452
rect 8364 9420 8393 9452
rect 8431 9420 8432 9452
rect 8432 9420 8465 9452
rect 8503 9420 8534 9452
rect 8534 9420 8537 9452
rect 8575 9420 8602 9452
rect 8602 9420 8609 9452
rect 8647 9420 8670 9452
rect 8670 9420 8681 9452
rect 8719 9420 8738 9452
rect 8738 9420 8753 9452
rect 8791 9420 8806 9452
rect 8806 9420 8825 9452
rect 8863 9420 8874 9452
rect 8874 9420 8897 9452
rect 8935 9420 8942 9452
rect 8942 9420 8969 9452
rect 9007 9420 9010 9452
rect 9010 9420 9041 9452
rect 9079 9420 9112 9452
rect 9112 9420 9113 9452
rect 9151 9420 9180 9452
rect 9180 9420 9185 9452
rect 9223 9420 9248 9452
rect 9248 9420 9257 9452
rect 9295 9420 9316 9452
rect 9316 9420 9329 9452
rect 9367 9420 9384 9452
rect 9384 9420 9401 9452
rect 9439 9420 9452 9452
rect 9452 9420 9473 9452
rect 9511 9420 9520 9452
rect 9520 9420 9545 9452
rect 9583 9420 9588 9452
rect 9588 9420 9617 9452
rect 9655 9420 9656 9452
rect 9656 9420 9689 9452
rect 9727 9420 9758 9452
rect 9758 9420 9761 9452
rect 9799 9420 9826 9452
rect 9826 9420 9833 9452
rect 9871 9420 9894 9452
rect 9894 9420 9905 9452
rect 9943 9420 9962 9452
rect 9962 9420 9977 9452
rect 10015 9420 10030 9452
rect 10030 9420 10049 9452
rect 10087 9420 10098 9452
rect 10098 9420 10121 9452
rect 10159 9420 10166 9452
rect 10166 9420 10193 9452
rect 10231 9420 10234 9452
rect 10234 9420 10265 9452
rect 10303 9420 10336 9452
rect 10336 9420 10337 9452
rect 10375 9420 10404 9452
rect 10404 9420 10409 9452
rect 10447 9420 10472 9452
rect 10472 9420 10481 9452
rect 10519 9420 10540 9452
rect 10540 9420 10553 9452
rect 10591 9420 10608 9452
rect 10608 9420 10625 9452
rect 10663 9420 10676 9452
rect 10676 9420 10697 9452
rect 10735 9420 10744 9452
rect 10744 9420 10769 9452
rect 10807 9420 10812 9452
rect 10812 9420 10841 9452
rect 10879 9420 10880 9452
rect 10880 9420 10913 9452
rect 10951 9420 10982 9452
rect 10982 9420 10985 9452
rect 11023 9420 11050 9452
rect 11050 9420 11057 9452
rect 11095 9420 11118 9452
rect 11118 9420 11129 9452
rect 11167 9420 11186 9452
rect 11186 9420 11201 9452
rect 11239 9420 11254 9452
rect 11254 9420 11273 9452
rect 11311 9420 11322 9452
rect 11322 9420 11345 9452
rect 11383 9420 11390 9452
rect 11390 9420 11417 9452
rect 11455 9420 11458 9452
rect 11458 9420 11489 9452
rect 11527 9420 11560 9452
rect 11560 9420 11561 9452
rect 11599 9420 11628 9452
rect 11628 9420 11633 9452
rect 11671 9420 11696 9452
rect 11696 9420 11705 9452
rect 11743 9420 11764 9452
rect 11764 9420 11777 9452
rect 11815 9420 11832 9452
rect 11832 9420 11849 9452
rect 11887 9420 11900 9452
rect 11900 9420 11921 9452
rect 11959 9420 11968 9452
rect 11968 9420 11993 9452
rect 12031 9420 12036 9452
rect 12036 9420 12065 9452
rect 12103 9420 12104 9452
rect 12104 9420 12137 9452
rect 12175 9420 12206 9452
rect 12206 9420 12209 9452
rect 12247 9420 12274 9452
rect 12274 9420 12281 9452
rect 12319 9420 12342 9452
rect 12342 9420 12353 9452
rect 12391 9420 12410 9452
rect 12410 9420 12425 9452
rect 12463 9420 12478 9452
rect 12478 9420 12497 9452
rect 12535 9420 12546 9452
rect 12546 9420 12569 9452
rect 12607 9420 12614 9452
rect 12614 9420 12641 9452
rect 14314 9420 14348 9452
rect 610 9418 644 9420
rect 2311 9418 2345 9420
rect 2383 9418 2417 9420
rect 2455 9418 2489 9420
rect 2527 9418 2561 9420
rect 2599 9418 2633 9420
rect 2671 9418 2705 9420
rect 2743 9418 2777 9420
rect 2815 9418 2849 9420
rect 2887 9418 2921 9420
rect 2959 9418 2993 9420
rect 3031 9418 3065 9420
rect 3103 9418 3137 9420
rect 3175 9418 3209 9420
rect 3247 9418 3281 9420
rect 3319 9418 3353 9420
rect 3391 9418 3425 9420
rect 3463 9418 3497 9420
rect 3535 9418 3569 9420
rect 3607 9418 3641 9420
rect 3679 9418 3713 9420
rect 3751 9418 3785 9420
rect 3823 9418 3857 9420
rect 3895 9418 3929 9420
rect 3967 9418 4001 9420
rect 4039 9418 4073 9420
rect 4111 9418 4145 9420
rect 4183 9418 4217 9420
rect 4255 9418 4289 9420
rect 4327 9418 4361 9420
rect 4399 9418 4433 9420
rect 4471 9418 4505 9420
rect 4543 9418 4577 9420
rect 4615 9418 4649 9420
rect 4687 9418 4721 9420
rect 4759 9418 4793 9420
rect 4831 9418 4865 9420
rect 4903 9418 4937 9420
rect 4975 9418 5009 9420
rect 5047 9418 5081 9420
rect 5119 9418 5153 9420
rect 5191 9418 5225 9420
rect 5263 9418 5297 9420
rect 5335 9418 5369 9420
rect 5407 9418 5441 9420
rect 5479 9418 5513 9420
rect 5551 9418 5585 9420
rect 5623 9418 5657 9420
rect 5695 9418 5729 9420
rect 5767 9418 5801 9420
rect 5839 9418 5873 9420
rect 5911 9418 5945 9420
rect 5983 9418 6017 9420
rect 6055 9418 6089 9420
rect 6127 9418 6161 9420
rect 6199 9418 6233 9420
rect 6271 9418 6305 9420
rect 6343 9418 6377 9420
rect 6415 9418 6449 9420
rect 6487 9418 6521 9420
rect 6559 9418 6593 9420
rect 6631 9418 6665 9420
rect 6703 9418 6737 9420
rect 6775 9418 6809 9420
rect 6847 9418 6881 9420
rect 6919 9418 6953 9420
rect 6991 9418 7025 9420
rect 7063 9418 7097 9420
rect 7135 9418 7169 9420
rect 7207 9418 7241 9420
rect 7279 9418 7313 9420
rect 7351 9418 7385 9420
rect 7423 9418 7457 9420
rect 7495 9418 7529 9420
rect 7567 9418 7601 9420
rect 7639 9418 7673 9420
rect 7711 9418 7745 9420
rect 7783 9418 7817 9420
rect 7855 9418 7889 9420
rect 7927 9418 7961 9420
rect 7999 9418 8033 9420
rect 8071 9418 8105 9420
rect 8143 9418 8177 9420
rect 8215 9418 8249 9420
rect 8287 9418 8321 9420
rect 8359 9418 8393 9420
rect 8431 9418 8465 9420
rect 8503 9418 8537 9420
rect 8575 9418 8609 9420
rect 8647 9418 8681 9420
rect 8719 9418 8753 9420
rect 8791 9418 8825 9420
rect 8863 9418 8897 9420
rect 8935 9418 8969 9420
rect 9007 9418 9041 9420
rect 9079 9418 9113 9420
rect 9151 9418 9185 9420
rect 9223 9418 9257 9420
rect 9295 9418 9329 9420
rect 9367 9418 9401 9420
rect 9439 9418 9473 9420
rect 9511 9418 9545 9420
rect 9583 9418 9617 9420
rect 9655 9418 9689 9420
rect 9727 9418 9761 9420
rect 9799 9418 9833 9420
rect 9871 9418 9905 9420
rect 9943 9418 9977 9420
rect 10015 9418 10049 9420
rect 10087 9418 10121 9420
rect 10159 9418 10193 9420
rect 10231 9418 10265 9420
rect 10303 9418 10337 9420
rect 10375 9418 10409 9420
rect 10447 9418 10481 9420
rect 10519 9418 10553 9420
rect 10591 9418 10625 9420
rect 10663 9418 10697 9420
rect 10735 9418 10769 9420
rect 10807 9418 10841 9420
rect 10879 9418 10913 9420
rect 10951 9418 10985 9420
rect 11023 9418 11057 9420
rect 11095 9418 11129 9420
rect 11167 9418 11201 9420
rect 11239 9418 11273 9420
rect 11311 9418 11345 9420
rect 11383 9418 11417 9420
rect 11455 9418 11489 9420
rect 11527 9418 11561 9420
rect 11599 9418 11633 9420
rect 11671 9418 11705 9420
rect 11743 9418 11777 9420
rect 11815 9418 11849 9420
rect 11887 9418 11921 9420
rect 11959 9418 11993 9420
rect 12031 9418 12065 9420
rect 12103 9418 12137 9420
rect 12175 9418 12209 9420
rect 12247 9418 12281 9420
rect 12319 9418 12353 9420
rect 12391 9418 12425 9420
rect 12463 9418 12497 9420
rect 12535 9418 12569 9420
rect 12607 9418 12641 9420
rect 14314 9418 14348 9420
rect 14614 9418 14648 9452
<< metal1 >>
rect 245 36534 14724 36574
rect 245 36500 320 36534
rect 354 36533 14724 36534
rect 354 36500 14614 36533
rect 245 36499 14614 36500
rect 14648 36499 14724 36533
rect 245 36498 14724 36499
rect 245 36464 556 36498
rect 590 36464 628 36498
rect 662 36464 700 36498
rect 734 36464 772 36498
rect 806 36464 844 36498
rect 878 36464 916 36498
rect 950 36464 988 36498
rect 1022 36464 1060 36498
rect 1094 36464 1132 36498
rect 1166 36464 1204 36498
rect 1238 36464 1276 36498
rect 1310 36464 1348 36498
rect 1382 36464 1420 36498
rect 1454 36464 1492 36498
rect 1526 36464 1564 36498
rect 1598 36464 1636 36498
rect 1670 36464 1708 36498
rect 1742 36464 1780 36498
rect 1814 36464 1852 36498
rect 1886 36464 1924 36498
rect 1958 36464 1996 36498
rect 2030 36464 2068 36498
rect 2102 36464 2140 36498
rect 2174 36464 2212 36498
rect 2246 36464 2284 36498
rect 2318 36464 2356 36498
rect 2390 36464 2428 36498
rect 2462 36464 2500 36498
rect 2534 36464 2572 36498
rect 2606 36464 2644 36498
rect 2678 36464 2716 36498
rect 2750 36464 2788 36498
rect 2822 36464 2860 36498
rect 2894 36464 2932 36498
rect 2966 36464 3004 36498
rect 3038 36464 3076 36498
rect 3110 36464 3148 36498
rect 3182 36464 3220 36498
rect 3254 36464 3292 36498
rect 3326 36464 3364 36498
rect 3398 36464 3436 36498
rect 3470 36464 3508 36498
rect 3542 36464 3580 36498
rect 3614 36464 3652 36498
rect 3686 36464 3724 36498
rect 3758 36464 3796 36498
rect 3830 36464 3868 36498
rect 3902 36464 3940 36498
rect 3974 36464 4012 36498
rect 4046 36464 4084 36498
rect 4118 36464 4156 36498
rect 4190 36464 4228 36498
rect 4262 36464 4300 36498
rect 4334 36464 4372 36498
rect 4406 36464 4444 36498
rect 4478 36464 4516 36498
rect 4550 36464 4588 36498
rect 4622 36464 4660 36498
rect 4694 36464 4732 36498
rect 4766 36464 4804 36498
rect 4838 36464 4876 36498
rect 4910 36464 4948 36498
rect 4982 36464 5020 36498
rect 5054 36464 5092 36498
rect 5126 36464 5164 36498
rect 5198 36464 5236 36498
rect 5270 36464 5308 36498
rect 5342 36464 5380 36498
rect 5414 36464 5452 36498
rect 5486 36464 5524 36498
rect 5558 36464 5596 36498
rect 5630 36464 5668 36498
rect 5702 36464 5740 36498
rect 5774 36464 5812 36498
rect 5846 36464 5884 36498
rect 5918 36464 5956 36498
rect 5990 36464 6028 36498
rect 6062 36464 6100 36498
rect 6134 36464 6172 36498
rect 6206 36464 6244 36498
rect 6278 36464 6316 36498
rect 6350 36464 6388 36498
rect 6422 36464 6460 36498
rect 6494 36464 6532 36498
rect 6566 36464 6604 36498
rect 6638 36464 6676 36498
rect 6710 36464 6748 36498
rect 6782 36464 6820 36498
rect 6854 36464 6892 36498
rect 6926 36464 6964 36498
rect 6998 36464 7036 36498
rect 7070 36464 7108 36498
rect 7142 36464 7180 36498
rect 7214 36464 7252 36498
rect 7286 36464 7324 36498
rect 7358 36464 7396 36498
rect 7430 36464 7468 36498
rect 7502 36464 7540 36498
rect 7574 36464 7612 36498
rect 7646 36464 7684 36498
rect 7718 36464 7756 36498
rect 7790 36464 7828 36498
rect 7862 36464 7900 36498
rect 7934 36464 7972 36498
rect 8006 36464 8044 36498
rect 8078 36464 8116 36498
rect 8150 36464 8188 36498
rect 8222 36464 8260 36498
rect 8294 36464 8332 36498
rect 8366 36464 8404 36498
rect 8438 36464 8476 36498
rect 8510 36464 8548 36498
rect 8582 36464 8620 36498
rect 8654 36464 8692 36498
rect 8726 36464 8764 36498
rect 8798 36464 8836 36498
rect 8870 36464 8908 36498
rect 8942 36464 8980 36498
rect 9014 36464 9052 36498
rect 9086 36464 9124 36498
rect 9158 36464 9196 36498
rect 9230 36464 9268 36498
rect 9302 36464 9340 36498
rect 9374 36464 9412 36498
rect 9446 36464 9484 36498
rect 9518 36464 9556 36498
rect 9590 36464 9628 36498
rect 9662 36464 9700 36498
rect 9734 36464 9772 36498
rect 9806 36464 9844 36498
rect 9878 36464 9916 36498
rect 9950 36464 9988 36498
rect 10022 36464 10060 36498
rect 10094 36464 10132 36498
rect 10166 36464 10204 36498
rect 10238 36464 10276 36498
rect 10310 36464 10348 36498
rect 10382 36464 10420 36498
rect 10454 36464 10492 36498
rect 10526 36464 10564 36498
rect 10598 36464 10636 36498
rect 10670 36464 10708 36498
rect 10742 36464 10780 36498
rect 10814 36464 10852 36498
rect 10886 36464 10924 36498
rect 10958 36464 10996 36498
rect 11030 36464 11068 36498
rect 11102 36464 11140 36498
rect 11174 36464 11212 36498
rect 11246 36464 11284 36498
rect 11318 36464 11356 36498
rect 11390 36464 11428 36498
rect 11462 36464 11500 36498
rect 11534 36464 11572 36498
rect 11606 36464 11644 36498
rect 11678 36464 11716 36498
rect 11750 36464 11788 36498
rect 11822 36464 11860 36498
rect 11894 36464 11932 36498
rect 11966 36464 12004 36498
rect 12038 36464 12076 36498
rect 12110 36464 12148 36498
rect 12182 36464 12220 36498
rect 12254 36464 12292 36498
rect 12326 36464 12364 36498
rect 12398 36464 12436 36498
rect 12470 36464 12508 36498
rect 12542 36464 12580 36498
rect 12614 36464 12652 36498
rect 12686 36464 12724 36498
rect 12758 36464 12796 36498
rect 12830 36464 12868 36498
rect 12902 36464 12940 36498
rect 12974 36464 13012 36498
rect 13046 36464 13084 36498
rect 13118 36464 13156 36498
rect 13190 36464 13228 36498
rect 13262 36464 13300 36498
rect 13334 36464 13372 36498
rect 13406 36464 13444 36498
rect 13478 36464 13516 36498
rect 13550 36464 13588 36498
rect 13622 36464 13660 36498
rect 13694 36464 13732 36498
rect 13766 36464 13804 36498
rect 13838 36464 13876 36498
rect 13910 36464 13948 36498
rect 13982 36464 14020 36498
rect 14054 36464 14092 36498
rect 14126 36464 14164 36498
rect 14198 36464 14236 36498
rect 14270 36464 14308 36498
rect 14342 36464 14380 36498
rect 14414 36464 14724 36498
rect 245 36462 14724 36464
rect 245 36428 320 36462
rect 354 36461 14724 36462
rect 354 36428 14614 36461
rect 245 36427 14614 36428
rect 14648 36427 14724 36461
rect 245 36389 14724 36427
rect 245 36265 430 36389
rect 245 36231 320 36265
rect 354 36231 430 36265
rect 245 36193 430 36231
rect 245 36159 320 36193
rect 354 36159 430 36193
rect 245 36121 430 36159
rect 245 36087 320 36121
rect 354 36087 430 36121
rect 245 36049 430 36087
rect 14539 36262 14724 36389
rect 14539 36228 14614 36262
rect 14648 36228 14724 36262
rect 14539 36190 14724 36228
rect 14539 36156 14614 36190
rect 14648 36156 14724 36190
rect 14539 36118 14724 36156
rect 14539 36084 14614 36118
rect 14648 36084 14724 36118
rect 245 36015 320 36049
rect 354 36015 430 36049
tri 850 36046 857 36053 se
rect 857 36046 14119 36053
tri 14119 36046 14126 36053 sw
rect 14539 36046 14724 36084
tri 823 36019 850 36046 se
rect 850 36019 14126 36046
rect 245 35977 430 36015
tri 816 36012 823 36019 se
rect 823 36012 14126 36019
tri 14126 36012 14160 36046 sw
rect 14539 36012 14614 36046
rect 14648 36012 14724 36046
tri 807 36003 816 36012 se
rect 816 36003 14160 36012
rect 245 35943 320 35977
rect 354 35943 430 35977
tri 773 35969 807 36003 se
rect 807 35969 1009 36003
rect 1043 35969 1081 36003
rect 1115 35969 1153 36003
rect 1187 35969 1225 36003
rect 1259 35969 1297 36003
rect 1331 35969 1369 36003
rect 1403 35969 1441 36003
rect 1475 35969 1513 36003
rect 1547 35969 1585 36003
rect 1619 35969 1657 36003
rect 1691 35969 1729 36003
rect 1763 35969 1801 36003
rect 1835 35969 1873 36003
rect 1907 35969 1945 36003
rect 1979 35969 2017 36003
rect 2051 35969 2089 36003
rect 2123 35969 2161 36003
rect 2195 35969 2233 36003
rect 2267 35969 2305 36003
rect 2339 35969 2377 36003
rect 2411 35969 2449 36003
rect 2483 35969 2521 36003
rect 2555 35969 2593 36003
rect 2627 35969 2665 36003
rect 2699 35969 2737 36003
rect 2771 35969 2809 36003
rect 2843 35969 2881 36003
rect 2915 35969 2953 36003
rect 2987 35969 3025 36003
rect 3059 35969 3097 36003
rect 3131 35969 3169 36003
rect 3203 35969 3241 36003
rect 3275 35969 3313 36003
rect 3347 35969 3385 36003
rect 3419 35969 3457 36003
rect 3491 35969 3529 36003
rect 3563 35969 3601 36003
rect 3635 35969 3673 36003
rect 3707 35969 3745 36003
rect 3779 35969 3817 36003
rect 3851 35969 3889 36003
rect 3923 35969 3961 36003
rect 3995 35969 4033 36003
rect 4067 35969 4105 36003
rect 4139 35969 4177 36003
rect 4211 35969 4249 36003
rect 4283 35969 4321 36003
rect 4355 35969 4393 36003
rect 4427 35969 4465 36003
rect 4499 35969 4537 36003
rect 4571 35969 4609 36003
rect 4643 35969 4681 36003
rect 4715 35969 4753 36003
rect 4787 35969 4825 36003
rect 4859 35969 4897 36003
rect 4931 35969 4969 36003
rect 5003 35969 5041 36003
rect 5075 35969 5113 36003
rect 5147 35969 5185 36003
rect 5219 35969 5257 36003
rect 5291 35969 5329 36003
rect 5363 35969 5401 36003
rect 5435 35969 5473 36003
rect 5507 35969 5545 36003
rect 5579 35969 5617 36003
rect 5651 35969 5689 36003
rect 5723 35969 5761 36003
rect 5795 35969 5833 36003
rect 5867 35969 5905 36003
rect 5939 35969 5977 36003
rect 6011 35969 6049 36003
rect 6083 35969 6121 36003
rect 6155 35969 6193 36003
rect 6227 35969 6265 36003
rect 6299 35969 6337 36003
rect 6371 35969 6409 36003
rect 6443 35969 6481 36003
rect 6515 35969 6553 36003
rect 6587 35969 6625 36003
rect 6659 35969 6697 36003
rect 6731 35969 6769 36003
rect 6803 35969 6841 36003
rect 6875 35969 6913 36003
rect 6947 35969 6985 36003
rect 7019 35969 7057 36003
rect 7091 35969 7129 36003
rect 7163 35969 7201 36003
rect 7235 35969 7273 36003
rect 7307 35969 7345 36003
rect 7379 35969 7417 36003
rect 7451 35969 7489 36003
rect 7523 35969 7561 36003
rect 7595 35969 7633 36003
rect 7667 35969 7705 36003
rect 7739 35969 7777 36003
rect 7811 35969 7849 36003
rect 7883 35969 7921 36003
rect 7955 35969 7993 36003
rect 8027 35969 8065 36003
rect 8099 35969 8137 36003
rect 8171 35969 8209 36003
rect 8243 35969 8281 36003
rect 8315 35969 8353 36003
rect 8387 35969 8425 36003
rect 8459 35969 8497 36003
rect 8531 35969 8569 36003
rect 8603 35969 8641 36003
rect 8675 35969 8713 36003
rect 8747 35969 8785 36003
rect 8819 35969 8857 36003
rect 8891 35969 8929 36003
rect 8963 35969 9001 36003
rect 9035 35969 9073 36003
rect 9107 35969 9145 36003
rect 9179 35969 9217 36003
rect 9251 35969 9289 36003
rect 9323 35969 9361 36003
rect 9395 35969 9433 36003
rect 9467 35969 9505 36003
rect 9539 35969 9577 36003
rect 9611 35969 9649 36003
rect 9683 35969 9721 36003
rect 9755 35969 9793 36003
rect 9827 35969 9865 36003
rect 9899 35969 9937 36003
rect 9971 35969 10009 36003
rect 10043 35969 10081 36003
rect 10115 35969 10153 36003
rect 10187 35969 10225 36003
rect 10259 35969 10297 36003
rect 10331 35969 10369 36003
rect 10403 35969 10441 36003
rect 10475 35969 10513 36003
rect 10547 35969 10585 36003
rect 10619 35969 10657 36003
rect 10691 35969 10729 36003
rect 10763 35969 10801 36003
rect 10835 35969 10873 36003
rect 10907 35969 10945 36003
rect 10979 35969 11017 36003
rect 11051 35969 11089 36003
rect 11123 35969 11161 36003
rect 11195 35969 11233 36003
rect 11267 35969 11305 36003
rect 11339 35969 11377 36003
rect 11411 35969 11449 36003
rect 11483 35969 11521 36003
rect 11555 35969 11593 36003
rect 11627 35969 11665 36003
rect 11699 35969 11737 36003
rect 11771 35969 11809 36003
rect 11843 35969 11881 36003
rect 11915 35969 11953 36003
rect 11987 35969 12025 36003
rect 12059 35969 12097 36003
rect 12131 35969 12169 36003
rect 12203 35969 12241 36003
rect 12275 35969 12313 36003
rect 12347 35969 12385 36003
rect 12419 35969 12457 36003
rect 12491 35969 12529 36003
rect 12563 35969 12601 36003
rect 12635 35969 12673 36003
rect 12707 35969 12745 36003
rect 12779 35969 12817 36003
rect 12851 35969 12889 36003
rect 12923 35969 12961 36003
rect 12995 35969 13033 36003
rect 13067 35969 13105 36003
rect 13139 35969 13177 36003
rect 13211 35969 13249 36003
rect 13283 35969 13321 36003
rect 13355 35969 13393 36003
rect 13427 35969 13465 36003
rect 13499 35969 13537 36003
rect 13571 35969 13609 36003
rect 13643 35969 13681 36003
rect 13715 35969 13753 36003
rect 13787 35969 13825 36003
rect 13859 35969 13897 36003
rect 13931 35969 13969 36003
rect 14003 35974 14160 36003
tri 14160 35974 14198 36012 sw
rect 14539 35974 14724 36012
rect 14003 35969 14198 35974
rect 245 35905 430 35943
rect 245 35871 320 35905
rect 354 35871 430 35905
rect 245 35833 430 35871
rect 245 35799 320 35833
rect 354 35799 430 35833
rect 245 35761 430 35799
rect 245 35727 320 35761
rect 354 35727 430 35761
rect 245 35689 430 35727
rect 245 35655 320 35689
rect 354 35655 430 35689
rect 245 35617 430 35655
rect 245 35583 320 35617
rect 354 35583 430 35617
rect 245 35545 430 35583
rect 245 35511 320 35545
rect 354 35511 430 35545
rect 245 35473 430 35511
rect 245 35439 320 35473
rect 354 35439 430 35473
rect 245 35401 430 35439
rect 245 35367 320 35401
rect 354 35367 430 35401
rect 245 35329 430 35367
rect 245 35295 320 35329
rect 354 35295 430 35329
rect 245 35257 430 35295
rect 245 35223 320 35257
rect 354 35223 430 35257
rect 245 35185 430 35223
rect 245 35151 320 35185
rect 354 35151 430 35185
rect 245 35113 430 35151
rect 245 35079 320 35113
rect 354 35079 430 35113
rect 245 35041 430 35079
rect 245 35007 320 35041
rect 354 35007 430 35041
rect 245 34969 430 35007
rect 245 34935 320 34969
rect 354 34935 430 34969
rect 245 34897 430 34935
rect 245 34863 320 34897
rect 354 34863 430 34897
rect 245 34825 430 34863
rect 245 34791 320 34825
rect 354 34791 430 34825
rect 245 34753 430 34791
rect 245 34719 320 34753
rect 354 34719 430 34753
rect 245 34681 430 34719
rect 245 34647 320 34681
rect 354 34647 430 34681
rect 245 34609 430 34647
rect 245 34575 320 34609
rect 354 34575 430 34609
rect 245 34537 430 34575
rect 245 34503 320 34537
rect 354 34503 430 34537
rect 245 34465 430 34503
rect 245 34431 320 34465
rect 354 34431 430 34465
rect 245 34393 430 34431
rect 245 34359 320 34393
rect 354 34359 430 34393
rect 245 34321 430 34359
rect 245 34287 320 34321
rect 354 34287 430 34321
rect 245 34249 430 34287
rect 245 34215 320 34249
rect 354 34215 430 34249
rect 245 34177 430 34215
rect 245 34143 320 34177
rect 354 34143 430 34177
rect 245 34105 430 34143
rect 245 34071 320 34105
rect 354 34071 430 34105
rect 245 34033 430 34071
rect 245 33999 320 34033
rect 354 33999 430 34033
rect 245 33961 430 33999
rect 245 33927 320 33961
rect 354 33927 430 33961
rect 245 33889 430 33927
rect 245 33855 320 33889
rect 354 33855 430 33889
rect 245 33817 430 33855
rect 245 33783 320 33817
rect 354 33783 430 33817
rect 245 33745 430 33783
rect 245 33711 320 33745
rect 354 33711 430 33745
rect 245 33673 430 33711
rect 245 33639 320 33673
rect 354 33639 430 33673
rect 245 33601 430 33639
rect 245 33567 320 33601
rect 354 33567 430 33601
rect 245 33529 430 33567
rect 245 33495 320 33529
rect 354 33495 430 33529
rect 245 33457 430 33495
rect 245 33423 320 33457
rect 354 33423 430 33457
rect 245 33385 430 33423
rect 245 33351 320 33385
rect 354 33351 430 33385
rect 245 33313 430 33351
rect 245 33279 320 33313
rect 354 33279 430 33313
rect 245 33241 430 33279
rect 245 33207 320 33241
rect 354 33207 430 33241
rect 245 33169 430 33207
rect 245 33135 320 33169
rect 354 33135 430 33169
rect 245 33097 430 33135
rect 245 33063 320 33097
rect 354 33063 430 33097
rect 245 33025 430 33063
rect 245 32991 320 33025
rect 354 32991 430 33025
rect 245 32953 430 32991
rect 245 32919 320 32953
rect 354 32919 430 32953
rect 245 32881 430 32919
rect 245 32847 320 32881
rect 354 32847 430 32881
rect 245 32809 430 32847
rect 245 32775 320 32809
rect 354 32775 430 32809
rect 245 32737 430 32775
rect 245 32703 320 32737
rect 354 32703 430 32737
rect 245 32665 430 32703
rect 245 32631 320 32665
rect 354 32631 430 32665
rect 245 32593 430 32631
rect 245 32559 320 32593
rect 354 32559 430 32593
rect 245 32521 430 32559
rect 245 32487 320 32521
rect 354 32487 430 32521
rect 245 32449 430 32487
rect 245 32415 320 32449
rect 354 32415 430 32449
rect 245 32377 430 32415
rect 245 32343 320 32377
rect 354 32343 430 32377
rect 245 32305 430 32343
rect 245 32271 320 32305
rect 354 32271 430 32305
rect 245 32233 430 32271
rect 245 32199 320 32233
rect 354 32199 430 32233
rect 245 32161 430 32199
rect 245 32127 320 32161
rect 354 32127 430 32161
rect 245 32089 430 32127
rect 245 32055 320 32089
rect 354 32055 430 32089
rect 245 32017 430 32055
rect 245 31983 320 32017
rect 354 31983 430 32017
rect 245 31945 430 31983
rect 245 31911 320 31945
rect 354 31911 430 31945
rect 245 31873 430 31911
rect 245 31839 320 31873
rect 354 31839 430 31873
rect 245 31801 430 31839
rect 245 31767 320 31801
rect 354 31767 430 31801
rect 245 31729 430 31767
rect 245 31695 320 31729
rect 354 31695 430 31729
rect 245 31657 430 31695
rect 245 31623 320 31657
rect 354 31623 430 31657
rect 245 31585 430 31623
rect 245 31551 320 31585
rect 354 31551 430 31585
rect 245 31513 430 31551
rect 245 31479 320 31513
rect 354 31479 430 31513
rect 245 31441 430 31479
rect 245 31407 320 31441
rect 354 31407 430 31441
rect 245 31369 430 31407
rect 245 31335 320 31369
rect 354 31335 430 31369
rect 245 31297 430 31335
rect 245 31263 320 31297
rect 354 31263 430 31297
rect 245 31225 430 31263
rect 245 31191 320 31225
rect 354 31191 430 31225
rect 245 31153 430 31191
rect 245 31119 320 31153
rect 354 31119 430 31153
rect 245 31081 430 31119
rect 245 31047 320 31081
rect 354 31047 430 31081
rect 245 31009 430 31047
rect 245 30975 320 31009
rect 354 30975 430 31009
rect 245 30937 430 30975
rect 245 30903 320 30937
rect 354 30903 430 30937
rect 245 30865 430 30903
rect 245 30831 320 30865
rect 354 30831 430 30865
rect 245 30793 430 30831
rect 245 30759 320 30793
rect 354 30759 430 30793
rect 245 30721 430 30759
rect 245 30687 320 30721
rect 354 30687 430 30721
rect 245 30649 430 30687
rect 245 30615 320 30649
rect 354 30615 430 30649
rect 245 30577 430 30615
rect 245 30543 320 30577
rect 354 30543 430 30577
rect 245 30505 430 30543
rect 245 30471 320 30505
rect 354 30471 430 30505
rect 245 30433 430 30471
rect 245 30399 320 30433
rect 354 30399 430 30433
rect 245 30361 430 30399
rect 245 30327 320 30361
rect 354 30327 430 30361
rect 245 30289 430 30327
rect 245 30255 320 30289
rect 354 30255 430 30289
rect 245 30217 430 30255
rect 245 30183 320 30217
rect 354 30183 430 30217
rect 245 30145 430 30183
rect 245 30111 320 30145
rect 354 30111 430 30145
rect 245 30073 430 30111
rect 245 30039 320 30073
rect 354 30039 430 30073
rect 245 30001 430 30039
rect 245 29967 320 30001
rect 354 29967 430 30001
rect 245 29929 430 29967
rect 245 29895 320 29929
rect 354 29895 430 29929
rect 245 29857 430 29895
rect 245 29823 320 29857
rect 354 29823 430 29857
rect 245 29785 430 29823
rect 245 29751 320 29785
rect 354 29751 430 29785
rect 245 29713 430 29751
rect 245 29679 320 29713
rect 354 29679 430 29713
rect 245 29641 430 29679
rect 245 29607 320 29641
rect 354 29607 430 29641
rect 245 29569 430 29607
rect 245 29535 320 29569
rect 354 29535 430 29569
rect 245 29497 430 29535
rect 245 29463 320 29497
rect 354 29463 430 29497
rect 245 29425 430 29463
rect 245 29391 320 29425
rect 354 29391 430 29425
rect 245 29353 430 29391
rect 245 29319 320 29353
rect 354 29319 430 29353
rect 245 29281 430 29319
rect 245 29247 320 29281
rect 354 29247 430 29281
rect 245 29209 430 29247
rect 245 29175 320 29209
rect 354 29175 430 29209
rect 245 29137 430 29175
rect 245 29103 320 29137
rect 354 29103 430 29137
rect 245 29065 430 29103
rect 245 29031 320 29065
rect 354 29031 430 29065
rect 245 28993 430 29031
rect 245 28959 320 28993
rect 354 28959 430 28993
rect 245 28921 430 28959
rect 245 28887 320 28921
rect 354 28887 430 28921
rect 245 28849 430 28887
rect 245 28815 320 28849
rect 354 28815 430 28849
rect 245 28777 430 28815
rect 245 28743 320 28777
rect 354 28743 430 28777
rect 245 28705 430 28743
rect 245 28671 320 28705
rect 354 28671 430 28705
rect 245 28633 430 28671
rect 245 28599 320 28633
rect 354 28599 430 28633
rect 245 28561 430 28599
rect 245 28527 320 28561
rect 354 28527 430 28561
rect 245 28489 430 28527
rect 245 28455 320 28489
rect 354 28455 430 28489
rect 245 28417 430 28455
rect 245 28383 320 28417
rect 354 28383 430 28417
rect 245 28345 430 28383
rect 245 28311 320 28345
rect 354 28311 430 28345
rect 245 28273 430 28311
rect 245 28239 320 28273
rect 354 28239 430 28273
rect 245 28201 430 28239
rect 245 28167 320 28201
rect 354 28167 430 28201
rect 245 28129 430 28167
rect 245 28095 320 28129
rect 354 28095 430 28129
rect 245 28057 430 28095
rect 245 28023 320 28057
rect 354 28023 430 28057
rect 245 27985 430 28023
rect 245 27951 320 27985
rect 354 27951 430 27985
rect 245 27913 430 27951
rect 245 27879 320 27913
rect 354 27879 430 27913
rect 245 27841 430 27879
rect 245 27807 320 27841
rect 354 27807 430 27841
rect 245 27769 430 27807
rect 245 27735 320 27769
rect 354 27735 430 27769
rect 245 27697 430 27735
rect 245 27663 320 27697
rect 354 27663 430 27697
rect 245 27625 430 27663
rect 245 27591 320 27625
rect 354 27591 430 27625
rect 245 27553 430 27591
rect 245 27519 320 27553
rect 354 27519 430 27553
rect 245 27481 430 27519
rect 245 27447 320 27481
rect 354 27447 430 27481
rect 245 27409 430 27447
rect 245 27375 320 27409
rect 354 27375 430 27409
rect 245 27337 430 27375
rect 245 27303 320 27337
rect 354 27303 430 27337
rect 245 27265 430 27303
rect 245 27231 320 27265
rect 354 27231 430 27265
rect 245 27193 430 27231
rect 245 27159 320 27193
rect 354 27159 430 27193
rect 245 27121 430 27159
rect 245 27087 320 27121
rect 354 27087 430 27121
rect 245 27049 430 27087
rect 245 27015 320 27049
rect 354 27015 430 27049
rect 245 26977 430 27015
rect 245 26943 320 26977
rect 354 26943 430 26977
rect 245 26905 430 26943
rect 245 26871 320 26905
rect 354 26871 430 26905
rect 245 26833 430 26871
rect 245 26799 320 26833
rect 354 26799 430 26833
rect 245 26761 430 26799
rect 245 26727 320 26761
rect 354 26727 430 26761
rect 245 26689 430 26727
rect 245 26655 320 26689
rect 354 26655 430 26689
rect 245 26617 430 26655
rect 245 26583 320 26617
rect 354 26583 430 26617
rect 245 26545 430 26583
rect 245 26511 320 26545
rect 354 26511 430 26545
rect 245 26473 430 26511
rect 245 26439 320 26473
rect 354 26439 430 26473
rect 245 26401 430 26439
rect 245 26367 320 26401
rect 354 26367 430 26401
rect 245 26329 430 26367
rect 245 26295 320 26329
rect 354 26295 430 26329
rect 245 26257 430 26295
rect 245 26223 320 26257
rect 354 26223 430 26257
rect 245 26185 430 26223
rect 245 26151 320 26185
rect 354 26151 430 26185
rect 245 26113 430 26151
rect 245 26079 320 26113
rect 354 26079 430 26113
rect 245 26041 430 26079
rect 245 26007 320 26041
rect 354 26007 430 26041
rect 245 25969 430 26007
rect 245 25935 320 25969
rect 354 25935 430 25969
rect 245 25897 430 25935
rect 245 25863 320 25897
rect 354 25863 430 25897
rect 245 25825 430 25863
rect 245 25791 320 25825
rect 354 25791 430 25825
rect 245 25753 430 25791
rect 245 25719 320 25753
rect 354 25719 430 25753
rect 245 25681 430 25719
rect 245 25647 320 25681
rect 354 25647 430 25681
rect 245 25609 430 25647
rect 245 25575 320 25609
rect 354 25575 430 25609
rect 245 25537 430 25575
rect 245 25503 320 25537
rect 354 25503 430 25537
rect 245 25465 430 25503
rect 245 25431 320 25465
rect 354 25431 430 25465
rect 245 25393 430 25431
rect 245 25359 320 25393
rect 354 25359 430 25393
rect 245 25321 430 25359
rect 245 25287 320 25321
rect 354 25287 430 25321
rect 245 25249 430 25287
rect 245 25215 320 25249
rect 354 25215 430 25249
rect 245 25177 430 25215
rect 245 25143 320 25177
rect 354 25143 430 25177
rect 245 25105 430 25143
rect 245 25071 320 25105
rect 354 25071 430 25105
rect 245 25033 430 25071
rect 245 24999 320 25033
rect 354 24999 430 25033
rect 245 24961 430 24999
rect 245 24927 320 24961
rect 354 24927 430 24961
rect 245 24889 430 24927
rect 245 24855 320 24889
rect 354 24855 430 24889
rect 245 24817 430 24855
rect 245 24783 320 24817
rect 354 24783 430 24817
rect 245 24745 430 24783
rect 245 24711 320 24745
rect 354 24711 430 24745
rect 245 24673 430 24711
rect 245 24639 320 24673
rect 354 24639 430 24673
rect 245 24601 430 24639
rect 245 24567 320 24601
rect 354 24567 430 24601
rect 245 24529 430 24567
rect 245 24495 320 24529
rect 354 24495 430 24529
rect 245 24457 430 24495
rect 245 24423 320 24457
rect 354 24423 430 24457
rect 245 24385 430 24423
rect 245 24351 320 24385
rect 354 24351 430 24385
rect 245 24313 430 24351
rect 245 24279 320 24313
rect 354 24279 430 24313
rect 245 24241 430 24279
rect 245 24207 320 24241
rect 354 24207 430 24241
rect 245 24169 430 24207
rect 245 24135 320 24169
rect 354 24135 430 24169
rect 245 24097 430 24135
rect 245 24063 320 24097
rect 354 24063 430 24097
rect 245 24025 430 24063
rect 245 23991 320 24025
rect 354 23991 430 24025
rect 245 23953 430 23991
rect 245 23919 320 23953
rect 354 23919 430 23953
rect 245 23881 430 23919
rect 245 23847 320 23881
rect 354 23847 430 23881
rect 245 23809 430 23847
rect 245 23775 320 23809
rect 354 23775 430 23809
rect 245 23737 430 23775
rect 245 23703 320 23737
rect 354 23703 430 23737
rect 245 23665 430 23703
rect 245 23631 320 23665
rect 354 23631 430 23665
rect 245 23593 430 23631
rect 245 23559 320 23593
rect 354 23559 430 23593
rect 245 23521 430 23559
rect 245 23487 320 23521
rect 354 23487 430 23521
rect 245 23449 430 23487
rect 245 23415 320 23449
rect 354 23415 430 23449
rect 245 23377 430 23415
rect 245 23343 320 23377
rect 354 23343 430 23377
rect 245 23305 430 23343
rect 245 23271 320 23305
rect 354 23271 430 23305
rect 245 23233 430 23271
rect 245 23199 320 23233
rect 354 23199 430 23233
rect 245 23161 430 23199
rect 245 23127 320 23161
rect 354 23127 430 23161
rect 245 23089 430 23127
rect 245 23055 320 23089
rect 354 23055 430 23089
rect 245 23017 430 23055
rect 245 22983 320 23017
rect 354 22983 430 23017
rect 245 22945 430 22983
rect 245 22911 320 22945
rect 354 22911 430 22945
rect 245 22873 430 22911
rect 245 22839 320 22873
rect 354 22839 430 22873
rect 245 22801 430 22839
rect 245 22767 320 22801
rect 354 22767 430 22801
rect 245 22729 430 22767
rect 245 22695 320 22729
rect 354 22695 430 22729
rect 245 22657 430 22695
rect 245 22623 320 22657
rect 354 22623 430 22657
rect 245 22585 430 22623
rect 245 22551 320 22585
rect 354 22551 430 22585
rect 245 22513 430 22551
rect 245 22479 320 22513
rect 354 22479 430 22513
rect 245 22441 430 22479
rect 245 22407 320 22441
rect 354 22407 430 22441
rect 245 22369 430 22407
rect 245 22335 320 22369
rect 354 22335 430 22369
rect 245 22297 430 22335
rect 245 22263 320 22297
rect 354 22263 430 22297
rect 245 22225 430 22263
rect 245 22191 320 22225
rect 354 22191 430 22225
rect 245 22153 430 22191
rect 245 22119 320 22153
rect 354 22119 430 22153
rect 245 22081 430 22119
rect 245 22047 320 22081
rect 354 22047 430 22081
rect 245 22009 430 22047
rect 245 21975 320 22009
rect 354 21975 430 22009
rect 245 21937 430 21975
rect 245 21903 320 21937
rect 354 21903 430 21937
rect 245 21865 430 21903
rect 245 21831 320 21865
rect 354 21831 430 21865
rect 245 21793 430 21831
rect 245 21759 320 21793
rect 354 21759 430 21793
rect 245 21721 430 21759
rect 245 21687 320 21721
rect 354 21687 430 21721
rect 245 21649 430 21687
rect 245 21615 320 21649
rect 354 21615 430 21649
rect 245 21577 430 21615
rect 245 21543 320 21577
rect 354 21543 430 21577
rect 245 21505 430 21543
rect 245 21471 320 21505
rect 354 21471 430 21505
rect 245 21433 430 21471
rect 245 21399 320 21433
rect 354 21399 430 21433
rect 245 21361 430 21399
rect 245 21327 320 21361
rect 354 21327 430 21361
rect 245 21289 430 21327
rect 245 21255 320 21289
rect 354 21255 430 21289
rect 245 21217 430 21255
rect 245 21183 320 21217
rect 354 21183 430 21217
rect 245 21145 430 21183
rect 245 21111 320 21145
rect 354 21111 430 21145
rect 245 21073 430 21111
rect 245 21039 320 21073
rect 354 21039 430 21073
rect 245 21001 430 21039
rect 245 20967 320 21001
rect 354 20967 430 21001
rect 245 20929 430 20967
rect 245 20895 320 20929
rect 354 20895 430 20929
rect 245 20857 430 20895
rect 245 20823 320 20857
rect 354 20823 430 20857
rect 245 20785 430 20823
rect 245 20751 320 20785
rect 354 20751 430 20785
rect 245 20713 430 20751
rect 245 20679 320 20713
rect 354 20679 430 20713
rect 245 20641 430 20679
rect 245 20607 320 20641
rect 354 20607 430 20641
rect 245 20569 430 20607
rect 245 20535 320 20569
rect 354 20535 430 20569
rect 245 20497 430 20535
rect 245 20463 320 20497
rect 354 20463 430 20497
rect 245 20425 430 20463
rect 245 20391 320 20425
rect 354 20391 430 20425
rect 245 20353 430 20391
rect 245 20319 320 20353
rect 354 20319 430 20353
rect 245 20281 430 20319
rect 245 20247 320 20281
rect 354 20247 430 20281
rect 245 20209 430 20247
rect 245 20175 320 20209
rect 354 20175 430 20209
rect 245 20137 430 20175
rect 245 20103 320 20137
rect 354 20103 430 20137
rect 245 20065 430 20103
rect 245 20031 320 20065
rect 354 20031 430 20065
rect 245 19993 430 20031
rect 245 19959 320 19993
rect 354 19959 430 19993
rect 245 19921 430 19959
rect 245 19887 320 19921
rect 354 19887 430 19921
rect 245 19849 430 19887
rect 245 19815 320 19849
rect 354 19815 430 19849
rect 245 19777 430 19815
rect 245 19743 320 19777
rect 354 19743 430 19777
rect 245 19705 430 19743
rect 245 19671 320 19705
rect 354 19671 430 19705
rect 245 19633 430 19671
rect 245 19599 320 19633
rect 354 19599 430 19633
rect 245 19561 430 19599
rect 245 19527 320 19561
rect 354 19527 430 19561
rect 245 19489 430 19527
rect 245 19455 320 19489
rect 354 19455 430 19489
rect 245 19417 430 19455
rect 245 19383 320 19417
rect 354 19383 430 19417
rect 245 19345 430 19383
rect 245 19311 320 19345
rect 354 19311 430 19345
rect 245 19273 430 19311
rect 245 19239 320 19273
rect 354 19239 430 19273
rect 245 19201 430 19239
rect 245 19167 320 19201
rect 354 19167 430 19201
rect 245 19129 430 19167
rect 245 19095 320 19129
rect 354 19095 430 19129
rect 245 19057 430 19095
rect 245 19023 320 19057
rect 354 19023 430 19057
rect 245 18985 430 19023
rect 245 18951 320 18985
rect 354 18951 430 18985
rect 245 18913 430 18951
rect 245 18879 320 18913
rect 354 18879 430 18913
rect 245 18841 430 18879
rect 245 18807 320 18841
rect 354 18807 430 18841
rect 245 18769 430 18807
rect 245 18735 320 18769
rect 354 18735 430 18769
rect 245 18697 430 18735
rect 245 18663 320 18697
rect 354 18663 430 18697
rect 245 18625 430 18663
rect 245 18591 320 18625
rect 354 18591 430 18625
rect 245 18553 430 18591
rect 245 18519 320 18553
rect 354 18519 430 18553
rect 245 18481 430 18519
rect 245 18447 320 18481
rect 354 18447 430 18481
rect 245 18409 430 18447
rect 245 18375 320 18409
rect 354 18375 430 18409
rect 245 18337 430 18375
rect 245 18303 320 18337
rect 354 18303 430 18337
rect 245 18265 430 18303
rect 245 18231 320 18265
rect 354 18231 430 18265
rect 245 18193 430 18231
rect 245 18159 320 18193
rect 354 18159 430 18193
rect 245 18121 430 18159
rect 245 18087 320 18121
rect 354 18087 430 18121
rect 245 18049 430 18087
rect 245 18015 320 18049
rect 354 18015 430 18049
rect 245 17977 430 18015
rect 245 17943 320 17977
rect 354 17943 430 17977
rect 245 17905 430 17943
rect 245 17871 320 17905
rect 354 17871 430 17905
rect 245 17833 430 17871
rect 245 17799 320 17833
rect 354 17799 430 17833
rect 245 17761 430 17799
rect 245 17727 320 17761
rect 354 17727 430 17761
rect 245 17689 430 17727
rect 245 17655 320 17689
rect 354 17655 430 17689
rect 245 17617 430 17655
rect 245 17583 320 17617
rect 354 17583 430 17617
rect 245 17545 430 17583
rect 245 17511 320 17545
rect 354 17511 430 17545
rect 245 17473 430 17511
rect 245 17439 320 17473
rect 354 17439 430 17473
rect 245 17401 430 17439
rect 245 17367 320 17401
rect 354 17367 430 17401
rect 245 17329 430 17367
rect 245 17295 320 17329
rect 354 17295 430 17329
rect 245 17257 430 17295
rect 245 17223 320 17257
rect 354 17223 430 17257
rect 245 17185 430 17223
rect 245 17151 320 17185
rect 354 17151 430 17185
rect 245 17113 430 17151
rect 245 17079 320 17113
rect 354 17079 430 17113
rect 245 17041 430 17079
rect 245 17007 320 17041
rect 354 17007 430 17041
rect 245 16969 430 17007
rect 245 16935 320 16969
rect 354 16935 430 16969
rect 245 16897 430 16935
rect 245 16863 320 16897
rect 354 16863 430 16897
rect 245 16825 430 16863
rect 245 16791 320 16825
rect 354 16791 430 16825
rect 245 16753 430 16791
rect 245 16719 320 16753
rect 354 16719 430 16753
rect 245 16681 430 16719
rect 245 16647 320 16681
rect 354 16647 430 16681
rect 245 16609 430 16647
rect 245 16575 320 16609
rect 354 16575 430 16609
rect 245 16537 430 16575
rect 245 16503 320 16537
rect 354 16503 430 16537
rect 245 16465 430 16503
rect 245 16431 320 16465
rect 354 16431 430 16465
rect 245 16393 430 16431
rect 245 16359 320 16393
rect 354 16359 430 16393
rect 245 16321 430 16359
rect 245 16287 320 16321
rect 354 16287 430 16321
rect 245 16249 430 16287
rect 245 16215 320 16249
rect 354 16215 430 16249
rect 245 16177 430 16215
rect 245 16143 320 16177
rect 354 16143 430 16177
rect 245 16105 430 16143
rect 245 16071 320 16105
rect 354 16071 430 16105
rect 245 16033 430 16071
rect 245 15999 320 16033
rect 354 15999 430 16033
rect 245 15961 430 15999
rect 245 15927 320 15961
rect 354 15927 430 15961
rect 245 15889 430 15927
rect 245 15855 320 15889
rect 354 15855 430 15889
rect 245 15817 430 15855
rect 245 15783 320 15817
rect 354 15783 430 15817
rect 245 15745 430 15783
rect 245 15711 320 15745
rect 354 15711 430 15745
rect 245 15673 430 15711
rect 245 15639 320 15673
rect 354 15639 430 15673
rect 245 15601 430 15639
rect 245 15567 320 15601
rect 354 15567 430 15601
rect 245 15529 430 15567
rect 245 15495 320 15529
rect 354 15495 430 15529
rect 245 15457 430 15495
rect 245 15423 320 15457
rect 354 15423 430 15457
rect 245 15385 430 15423
rect 245 15351 320 15385
rect 354 15351 430 15385
rect 245 15313 430 15351
rect 245 15279 320 15313
rect 354 15279 430 15313
rect 245 15241 430 15279
rect 245 15207 320 15241
rect 354 15207 430 15241
rect 245 15169 430 15207
rect 245 15135 320 15169
rect 354 15135 430 15169
rect 245 15097 430 15135
rect 245 15063 320 15097
rect 354 15063 430 15097
rect 245 15025 430 15063
rect 245 14991 320 15025
rect 354 14991 430 15025
rect 245 14953 430 14991
rect 245 14919 320 14953
rect 354 14919 430 14953
rect 245 14881 430 14919
rect 245 14847 320 14881
rect 354 14847 430 14881
rect 245 14809 430 14847
rect 245 14775 320 14809
rect 354 14775 430 14809
rect 245 14737 430 14775
rect 245 14703 320 14737
rect 354 14703 430 14737
rect 245 14665 430 14703
rect 245 14631 320 14665
rect 354 14631 430 14665
rect 245 14593 430 14631
rect 245 14559 320 14593
rect 354 14559 430 14593
rect 245 14521 430 14559
rect 245 14487 320 14521
rect 354 14487 430 14521
rect 245 14449 430 14487
rect 245 14415 320 14449
rect 354 14415 430 14449
rect 245 14377 430 14415
rect 245 14343 320 14377
rect 354 14343 430 14377
rect 245 14305 430 14343
rect 245 14271 320 14305
rect 354 14271 430 14305
rect 245 14233 430 14271
rect 245 14199 320 14233
rect 354 14199 430 14233
rect 245 14161 430 14199
rect 245 14127 320 14161
rect 354 14127 430 14161
rect 245 14089 430 14127
rect 245 14055 320 14089
rect 354 14055 430 14089
rect 245 14017 430 14055
rect 245 13983 320 14017
rect 354 13983 430 14017
rect 245 13945 430 13983
rect 245 13911 320 13945
rect 354 13911 430 13945
rect 245 13873 430 13911
rect 245 13839 320 13873
rect 354 13839 430 13873
rect 245 13801 430 13839
rect 245 13767 320 13801
rect 354 13767 430 13801
rect 245 13729 430 13767
rect 245 13695 320 13729
rect 354 13695 430 13729
rect 245 13657 430 13695
rect 245 13623 320 13657
rect 354 13623 430 13657
rect 245 13585 430 13623
rect 245 13551 320 13585
rect 354 13551 430 13585
rect 245 13513 430 13551
rect 245 13479 320 13513
rect 354 13479 430 13513
rect 245 13441 430 13479
rect 245 13407 320 13441
rect 354 13407 430 13441
rect 245 13369 430 13407
rect 245 13335 320 13369
rect 354 13335 430 13369
rect 245 13297 430 13335
rect 245 13263 320 13297
rect 354 13263 430 13297
rect 245 13225 430 13263
rect 245 13191 320 13225
rect 354 13191 430 13225
rect 245 13153 430 13191
rect 245 13119 320 13153
rect 354 13119 430 13153
rect 245 13081 430 13119
rect 245 13047 320 13081
rect 354 13047 430 13081
rect 245 13009 430 13047
rect 245 12975 320 13009
rect 354 12975 430 13009
rect 245 12937 430 12975
rect 245 12903 320 12937
rect 354 12903 430 12937
rect 245 12865 430 12903
rect 245 12831 320 12865
rect 354 12831 430 12865
rect 245 12793 430 12831
rect 245 12759 320 12793
rect 354 12759 430 12793
rect 245 12721 430 12759
rect 245 12687 320 12721
rect 354 12687 430 12721
rect 245 12649 430 12687
rect 245 12615 320 12649
rect 354 12615 430 12649
rect 245 12577 430 12615
rect 245 12543 320 12577
rect 354 12543 430 12577
rect 245 12505 430 12543
rect 245 12471 320 12505
rect 354 12471 430 12505
rect 245 12433 430 12471
rect 245 12399 320 12433
rect 354 12399 430 12433
rect 245 12361 430 12399
rect 245 12327 320 12361
rect 354 12327 430 12361
rect 245 12289 430 12327
rect 245 12255 320 12289
rect 354 12255 430 12289
rect 245 12217 430 12255
rect 245 12183 320 12217
rect 354 12183 430 12217
rect 245 12145 430 12183
rect 245 12111 320 12145
rect 354 12111 430 12145
rect 245 12073 430 12111
rect 245 12039 320 12073
rect 354 12039 430 12073
rect 245 12001 430 12039
rect 245 11967 320 12001
rect 354 11967 430 12001
rect 245 11929 430 11967
rect 245 11895 320 11929
rect 354 11895 430 11929
rect 245 11857 430 11895
rect 245 11823 320 11857
rect 354 11823 430 11857
rect 245 11785 430 11823
rect 245 11751 320 11785
rect 354 11751 430 11785
rect 245 11713 430 11751
rect 245 11679 320 11713
rect 354 11679 430 11713
rect 245 11641 430 11679
rect 245 11607 320 11641
rect 354 11607 430 11641
rect 245 11569 430 11607
rect 245 11535 320 11569
rect 354 11535 430 11569
rect 245 11497 430 11535
rect 245 11463 320 11497
rect 354 11463 430 11497
rect 245 11425 430 11463
rect 245 11391 320 11425
rect 354 11391 430 11425
rect 245 11353 430 11391
rect 245 11319 320 11353
rect 354 11319 430 11353
rect 245 11281 430 11319
rect 245 11247 320 11281
rect 354 11247 430 11281
rect 245 11209 430 11247
rect 245 11175 320 11209
rect 354 11175 430 11209
rect 245 11137 430 11175
rect 245 11103 320 11137
rect 354 11103 430 11137
rect 245 11065 430 11103
rect 245 11031 320 11065
rect 354 11031 430 11065
rect 245 10993 430 11031
rect 245 10959 320 10993
rect 354 10959 430 10993
rect 245 10921 430 10959
rect 245 10887 320 10921
rect 354 10887 430 10921
rect 245 10849 430 10887
rect 245 10815 320 10849
rect 354 10815 430 10849
rect 245 10777 430 10815
rect 245 10743 320 10777
rect 354 10743 430 10777
rect 245 10705 430 10743
rect 245 10671 320 10705
rect 354 10671 430 10705
rect 245 10633 430 10671
rect 245 10599 320 10633
rect 354 10599 430 10633
rect 245 10561 430 10599
rect 245 10527 320 10561
rect 354 10527 430 10561
rect 245 10489 430 10527
rect 245 10455 320 10489
rect 354 10455 430 10489
rect 245 10417 430 10455
rect 245 10383 320 10417
rect 354 10383 430 10417
rect 245 10345 430 10383
rect 245 10311 320 10345
rect 354 10311 430 10345
rect 245 10273 430 10311
rect 245 10239 320 10273
rect 354 10239 430 10273
rect 245 10201 430 10239
rect 245 10167 320 10201
rect 354 10167 430 10201
rect 245 10129 430 10167
rect 245 10095 320 10129
rect 354 10095 430 10129
rect 245 10057 430 10095
rect 245 10023 320 10057
rect 354 10023 430 10057
rect 245 9985 430 10023
rect 245 9951 320 9985
rect 354 9951 430 9985
rect 245 9913 430 9951
tri 757 35953 773 35969 se
rect 773 35953 14198 35969
tri 14198 35953 14219 35974 sw
rect 757 35933 14219 35953
rect 757 35911 886 35933
rect 757 35877 814 35911
rect 848 35902 886 35911
tri 886 35902 917 35933 nw
tri 14059 35902 14090 35933 ne
rect 14090 35902 14219 35933
rect 848 35877 877 35902
tri 877 35893 886 35902 nw
tri 14090 35893 14099 35902 ne
rect 757 35839 877 35877
rect 757 35805 814 35839
rect 848 35805 877 35839
rect 757 35767 877 35805
rect 757 35733 814 35767
rect 848 35733 877 35767
rect 757 35695 877 35733
rect 757 35661 814 35695
rect 848 35661 877 35695
rect 757 35623 877 35661
rect 757 35589 814 35623
rect 848 35589 877 35623
rect 757 35551 877 35589
rect 757 35517 814 35551
rect 848 35517 877 35551
rect 757 35479 877 35517
rect 757 35445 814 35479
rect 848 35445 877 35479
rect 757 35407 877 35445
rect 757 35373 814 35407
rect 848 35373 877 35407
rect 757 35335 877 35373
rect 757 35301 814 35335
rect 848 35301 877 35335
rect 757 35263 877 35301
rect 757 35229 814 35263
rect 848 35229 877 35263
rect 757 35191 877 35229
rect 757 35157 814 35191
rect 848 35157 877 35191
rect 757 35119 877 35157
rect 757 35085 814 35119
rect 848 35085 877 35119
rect 757 35047 877 35085
rect 757 35013 814 35047
rect 848 35013 877 35047
rect 757 34975 877 35013
rect 757 34941 814 34975
rect 848 34941 877 34975
rect 757 34903 877 34941
rect 757 34869 814 34903
rect 848 34869 877 34903
rect 757 34831 877 34869
rect 757 34797 814 34831
rect 848 34797 877 34831
rect 757 34759 877 34797
rect 757 34725 814 34759
rect 848 34725 877 34759
rect 757 34687 877 34725
rect 757 34653 814 34687
rect 848 34653 877 34687
rect 14099 35832 14219 35902
rect 14099 35798 14120 35832
rect 14154 35798 14219 35832
rect 14099 35760 14219 35798
rect 14099 35726 14120 35760
rect 14154 35726 14219 35760
rect 14099 35688 14219 35726
rect 14099 35654 14120 35688
rect 14154 35654 14219 35688
rect 14099 35616 14219 35654
rect 14099 35582 14120 35616
rect 14154 35582 14219 35616
rect 14099 35544 14219 35582
rect 14099 35510 14120 35544
rect 14154 35510 14219 35544
rect 14099 35472 14219 35510
rect 14099 35438 14120 35472
rect 14154 35438 14219 35472
rect 14099 35400 14219 35438
rect 14099 35366 14120 35400
rect 14154 35366 14219 35400
rect 14099 35328 14219 35366
rect 14099 35294 14120 35328
rect 14154 35294 14219 35328
rect 14099 35256 14219 35294
rect 14099 35222 14120 35256
rect 14154 35222 14219 35256
rect 14099 35184 14219 35222
rect 14099 35150 14120 35184
rect 14154 35150 14219 35184
rect 14099 35112 14219 35150
rect 14099 35078 14120 35112
rect 14154 35078 14219 35112
rect 14099 35040 14219 35078
rect 14099 35006 14120 35040
rect 14154 35006 14219 35040
rect 14099 34968 14219 35006
rect 14099 34934 14120 34968
rect 14154 34934 14219 34968
rect 14099 34896 14219 34934
rect 14099 34862 14120 34896
rect 14154 34862 14219 34896
rect 14099 34824 14219 34862
rect 14099 34790 14120 34824
rect 14154 34790 14219 34824
rect 14099 34752 14219 34790
rect 14099 34718 14120 34752
rect 14154 34718 14219 34752
rect 757 34615 877 34653
rect 757 34581 814 34615
rect 848 34581 877 34615
rect 757 34543 877 34581
rect 757 34509 814 34543
rect 848 34509 877 34543
rect 757 34471 877 34509
rect 757 34437 814 34471
rect 848 34437 877 34471
rect 757 34399 877 34437
rect 757 34365 814 34399
rect 848 34365 877 34399
rect 757 34327 877 34365
rect 757 34293 814 34327
rect 848 34293 877 34327
rect 757 34255 877 34293
rect 757 34221 814 34255
rect 848 34221 877 34255
rect 757 34183 877 34221
rect 757 34149 814 34183
rect 848 34149 877 34183
rect 757 34111 877 34149
rect 757 34077 814 34111
rect 848 34077 877 34111
rect 757 34039 877 34077
rect 757 34005 814 34039
rect 848 34005 877 34039
rect 757 33967 877 34005
rect 757 33933 814 33967
rect 848 33933 877 33967
rect 757 33895 877 33933
rect 757 33861 814 33895
rect 848 33861 877 33895
rect 757 33823 877 33861
rect 757 33789 814 33823
rect 848 33789 877 33823
rect 757 33751 877 33789
rect 757 33717 814 33751
rect 848 33717 877 33751
rect 757 33679 877 33717
rect 757 33645 814 33679
rect 848 33645 877 33679
rect 757 33607 877 33645
rect 757 33573 814 33607
rect 848 33573 877 33607
rect 757 33535 877 33573
rect 757 33501 814 33535
rect 848 33501 877 33535
rect 757 33463 877 33501
rect 757 33429 814 33463
rect 848 33429 877 33463
rect 757 33391 877 33429
rect 757 33357 814 33391
rect 848 33357 877 33391
rect 757 33319 877 33357
rect 757 33285 814 33319
rect 848 33285 877 33319
rect 757 33247 877 33285
rect 757 33213 814 33247
rect 848 33213 877 33247
rect 757 33175 877 33213
rect 757 33141 814 33175
rect 848 33141 877 33175
rect 757 33103 877 33141
rect 757 33069 814 33103
rect 848 33069 877 33103
rect 757 33031 877 33069
rect 757 32997 814 33031
rect 848 32997 877 33031
rect 757 32959 877 32997
rect 757 32925 814 32959
rect 848 32925 877 32959
rect 757 32887 877 32925
rect 757 32853 814 32887
rect 848 32853 877 32887
rect 757 32815 877 32853
rect 757 32781 814 32815
rect 848 32781 877 32815
rect 757 32743 877 32781
rect 757 32709 814 32743
rect 848 32709 877 32743
rect 757 32671 877 32709
rect 757 32637 814 32671
rect 848 32637 877 32671
rect 757 32599 877 32637
rect 757 32565 814 32599
rect 848 32565 877 32599
rect 757 32527 877 32565
rect 757 32493 814 32527
rect 848 32493 877 32527
rect 757 32455 877 32493
rect 757 32421 814 32455
rect 848 32421 877 32455
rect 757 32383 877 32421
rect 757 32349 814 32383
rect 848 32349 877 32383
rect 757 32311 877 32349
rect 757 32277 814 32311
rect 848 32277 877 32311
rect 757 32239 877 32277
rect 757 32205 814 32239
rect 848 32205 877 32239
rect 757 32167 877 32205
rect 757 32133 814 32167
rect 848 32133 877 32167
rect 757 32095 877 32133
rect 757 32061 814 32095
rect 848 32061 877 32095
rect 757 32023 877 32061
rect 757 31989 814 32023
rect 848 31989 877 32023
rect 757 31951 877 31989
rect 757 31917 814 31951
rect 848 31917 877 31951
rect 757 31879 877 31917
rect 757 31845 814 31879
rect 848 31845 877 31879
rect 757 31807 877 31845
rect 757 31773 814 31807
rect 848 31773 877 31807
rect 757 31735 877 31773
rect 757 31701 814 31735
rect 848 31701 877 31735
rect 757 31663 877 31701
rect 757 31629 814 31663
rect 848 31629 877 31663
rect 757 31591 877 31629
rect 757 31557 814 31591
rect 848 31557 877 31591
rect 757 31519 877 31557
rect 757 31485 814 31519
rect 848 31485 877 31519
rect 757 31447 877 31485
rect 757 31413 814 31447
rect 848 31413 877 31447
rect 757 31375 877 31413
rect 757 31341 814 31375
rect 848 31341 877 31375
rect 757 31303 877 31341
rect 757 31269 814 31303
rect 848 31269 877 31303
rect 757 31231 877 31269
rect 757 31197 814 31231
rect 848 31197 877 31231
rect 757 31159 877 31197
rect 757 31125 814 31159
rect 848 31125 877 31159
rect 757 31087 877 31125
rect 757 31053 814 31087
rect 848 31053 877 31087
rect 757 31015 877 31053
rect 757 30981 814 31015
rect 848 30981 877 31015
rect 757 30943 877 30981
rect 757 30909 814 30943
rect 848 30909 877 30943
rect 757 30871 877 30909
rect 757 30837 814 30871
rect 848 30837 877 30871
rect 757 30799 877 30837
rect 757 30765 814 30799
rect 848 30765 877 30799
rect 757 30727 877 30765
rect 757 30693 814 30727
rect 848 30693 877 30727
rect 757 30655 877 30693
rect 757 30621 814 30655
rect 848 30621 877 30655
rect 757 30583 877 30621
rect 757 30549 814 30583
rect 848 30549 877 30583
rect 757 30511 877 30549
rect 757 30477 814 30511
rect 848 30477 877 30511
rect 757 30439 877 30477
rect 757 30405 814 30439
rect 848 30405 877 30439
rect 757 30367 877 30405
rect 757 30333 814 30367
rect 848 30333 877 30367
rect 757 30295 877 30333
rect 757 30261 814 30295
rect 848 30261 877 30295
rect 757 30223 877 30261
rect 757 30189 814 30223
rect 848 30189 877 30223
rect 757 30151 877 30189
rect 757 30117 814 30151
rect 848 30117 877 30151
rect 757 30079 877 30117
rect 757 30045 814 30079
rect 848 30045 877 30079
rect 757 30007 877 30045
rect 757 29973 814 30007
rect 848 29973 877 30007
rect 757 29935 877 29973
rect 757 29901 814 29935
rect 848 29901 877 29935
rect 757 29863 877 29901
rect 757 29829 814 29863
rect 848 29829 877 29863
rect 757 29791 877 29829
rect 757 29757 814 29791
rect 848 29757 877 29791
rect 757 29719 877 29757
rect 757 29685 814 29719
rect 848 29685 877 29719
rect 757 29647 877 29685
rect 757 29613 814 29647
rect 848 29613 877 29647
rect 757 29575 877 29613
rect 757 29541 814 29575
rect 848 29541 877 29575
rect 757 29503 877 29541
rect 757 29469 814 29503
rect 848 29469 877 29503
rect 757 29431 877 29469
rect 757 29397 814 29431
rect 848 29397 877 29431
rect 757 29359 877 29397
rect 757 29325 814 29359
rect 848 29325 877 29359
rect 757 29287 877 29325
rect 757 29253 814 29287
rect 848 29253 877 29287
rect 757 29215 877 29253
rect 757 29181 814 29215
rect 848 29181 877 29215
rect 757 29143 877 29181
rect 757 29109 814 29143
rect 848 29109 877 29143
rect 757 29071 877 29109
rect 757 29037 814 29071
rect 848 29037 877 29071
rect 757 28999 877 29037
rect 757 28965 814 28999
rect 848 28965 877 28999
rect 757 28927 877 28965
rect 757 28893 814 28927
rect 848 28893 877 28927
rect 757 28855 877 28893
rect 757 28821 814 28855
rect 848 28821 877 28855
rect 757 28783 877 28821
rect 757 28749 814 28783
rect 848 28749 877 28783
rect 757 28711 877 28749
rect 757 28677 814 28711
rect 848 28677 877 28711
rect 757 28639 877 28677
rect 757 28605 814 28639
rect 848 28605 877 28639
rect 757 28567 877 28605
rect 757 28533 814 28567
rect 848 28533 877 28567
rect 757 28495 877 28533
rect 757 28461 814 28495
rect 848 28461 877 28495
rect 757 28423 877 28461
rect 757 28389 814 28423
rect 848 28389 877 28423
rect 757 28351 877 28389
rect 757 28317 814 28351
rect 848 28317 877 28351
rect 757 28279 877 28317
rect 757 28245 814 28279
rect 848 28245 877 28279
rect 757 28207 877 28245
rect 757 28173 814 28207
rect 848 28173 877 28207
rect 757 28135 877 28173
rect 757 28101 814 28135
rect 848 28101 877 28135
rect 757 28063 877 28101
rect 757 28029 814 28063
rect 848 28029 877 28063
rect 757 27991 877 28029
rect 757 27957 814 27991
rect 848 27957 877 27991
rect 757 27919 877 27957
rect 757 27885 814 27919
rect 848 27885 877 27919
rect 757 27847 877 27885
rect 757 27813 814 27847
rect 848 27813 877 27847
rect 757 27775 877 27813
rect 757 27741 814 27775
rect 848 27741 877 27775
rect 757 27703 877 27741
rect 757 27669 814 27703
rect 848 27669 877 27703
rect 757 27631 877 27669
rect 757 27597 814 27631
rect 848 27597 877 27631
rect 757 27559 877 27597
rect 757 27525 814 27559
rect 848 27525 877 27559
rect 757 27487 877 27525
rect 757 27453 814 27487
rect 848 27453 877 27487
rect 757 27415 877 27453
rect 757 27381 814 27415
rect 848 27381 877 27415
rect 757 27343 877 27381
rect 757 27309 814 27343
rect 848 27309 877 27343
rect 757 27271 877 27309
rect 757 27237 814 27271
rect 848 27237 877 27271
rect 757 27199 877 27237
rect 757 27165 814 27199
rect 848 27165 877 27199
rect 757 27127 877 27165
rect 757 27093 814 27127
rect 848 27093 877 27127
rect 757 27055 877 27093
rect 757 27021 814 27055
rect 848 27021 877 27055
rect 757 26983 877 27021
rect 757 26949 814 26983
rect 848 26949 877 26983
rect 757 26911 877 26949
rect 757 26877 814 26911
rect 848 26877 877 26911
rect 757 26839 877 26877
rect 757 26805 814 26839
rect 848 26805 877 26839
rect 757 26767 877 26805
rect 757 26733 814 26767
rect 848 26733 877 26767
rect 757 26695 877 26733
rect 757 26661 814 26695
rect 848 26661 877 26695
rect 757 26623 877 26661
rect 757 26589 814 26623
rect 848 26589 877 26623
rect 757 26551 877 26589
rect 757 26517 814 26551
rect 848 26517 877 26551
rect 757 26479 877 26517
rect 757 26445 814 26479
rect 848 26445 877 26479
rect 757 26407 877 26445
rect 757 26373 814 26407
rect 848 26373 877 26407
rect 757 26335 877 26373
rect 757 26301 814 26335
rect 848 26301 877 26335
rect 757 26263 877 26301
rect 757 26229 814 26263
rect 848 26229 877 26263
rect 757 26191 877 26229
rect 757 26157 814 26191
rect 848 26157 877 26191
rect 757 26119 877 26157
rect 757 26085 814 26119
rect 848 26085 877 26119
rect 757 26047 877 26085
rect 757 26013 814 26047
rect 848 26013 877 26047
rect 757 25975 877 26013
rect 757 25941 814 25975
rect 848 25941 877 25975
rect 757 25903 877 25941
rect 757 25869 814 25903
rect 848 25869 877 25903
rect 757 25831 877 25869
rect 757 25797 814 25831
rect 848 25797 877 25831
rect 757 25759 877 25797
rect 757 25725 814 25759
rect 848 25725 877 25759
rect 757 25687 877 25725
rect 757 25653 814 25687
rect 848 25653 877 25687
rect 757 25615 877 25653
rect 757 25581 814 25615
rect 848 25581 877 25615
rect 757 25543 877 25581
rect 757 25509 814 25543
rect 848 25509 877 25543
rect 757 25471 877 25509
rect 757 25437 814 25471
rect 848 25437 877 25471
rect 757 25399 877 25437
rect 757 25365 814 25399
rect 848 25365 877 25399
rect 757 25327 877 25365
rect 757 25293 814 25327
rect 848 25293 877 25327
rect 757 25255 877 25293
rect 757 25221 814 25255
rect 848 25221 877 25255
rect 757 25183 877 25221
rect 757 25149 814 25183
rect 848 25149 877 25183
rect 757 25111 877 25149
rect 757 25077 814 25111
rect 848 25077 877 25111
rect 757 25039 877 25077
rect 757 25005 814 25039
rect 848 25005 877 25039
rect 757 24967 877 25005
rect 757 24933 814 24967
rect 848 24933 877 24967
rect 757 24895 877 24933
rect 757 24861 814 24895
rect 848 24861 877 24895
rect 757 24823 877 24861
rect 757 24789 814 24823
rect 848 24789 877 24823
rect 757 24751 877 24789
rect 757 24717 814 24751
rect 848 24717 877 24751
rect 757 24679 877 24717
rect 757 24645 814 24679
rect 848 24645 877 24679
rect 757 24607 877 24645
rect 757 24573 814 24607
rect 848 24573 877 24607
rect 757 24535 877 24573
rect 757 24501 814 24535
rect 848 24501 877 24535
rect 757 24463 877 24501
rect 757 24429 814 24463
rect 848 24429 877 24463
rect 757 24391 877 24429
rect 757 24357 814 24391
rect 848 24357 877 24391
rect 757 24319 877 24357
rect 757 24285 814 24319
rect 848 24285 877 24319
rect 757 24247 877 24285
rect 757 24213 814 24247
rect 848 24213 877 24247
rect 757 24175 877 24213
rect 757 24141 814 24175
rect 848 24141 877 24175
rect 757 24103 877 24141
rect 757 24069 814 24103
rect 848 24069 877 24103
rect 757 24031 877 24069
rect 757 23997 814 24031
rect 848 23997 877 24031
rect 757 23959 877 23997
rect 757 23925 814 23959
rect 848 23925 877 23959
rect 757 23887 877 23925
rect 757 23853 814 23887
rect 848 23853 877 23887
rect 757 23815 877 23853
rect 757 23781 814 23815
rect 848 23781 877 23815
rect 757 23743 877 23781
rect 757 23709 814 23743
rect 848 23709 877 23743
rect 757 23671 877 23709
rect 757 23637 814 23671
rect 848 23637 877 23671
rect 757 23599 877 23637
rect 757 23565 814 23599
rect 848 23565 877 23599
rect 757 23527 877 23565
rect 757 23493 814 23527
rect 848 23493 877 23527
rect 757 23455 877 23493
rect 757 23421 814 23455
rect 848 23421 877 23455
rect 757 23383 877 23421
rect 757 23349 814 23383
rect 848 23349 877 23383
rect 757 23311 877 23349
rect 757 23277 814 23311
rect 848 23277 877 23311
rect 757 23239 877 23277
rect 757 23205 814 23239
rect 848 23205 877 23239
rect 757 23167 877 23205
rect 757 23133 814 23167
rect 848 23133 877 23167
rect 757 23095 877 23133
rect 757 23061 814 23095
rect 848 23061 877 23095
rect 757 23023 877 23061
rect 757 22989 814 23023
rect 848 22989 877 23023
rect 757 22951 877 22989
rect 757 22917 814 22951
rect 848 22917 877 22951
rect 757 22879 877 22917
rect 757 22845 814 22879
rect 848 22845 877 22879
rect 757 22807 877 22845
rect 757 22773 814 22807
rect 848 22773 877 22807
rect 757 22735 877 22773
rect 757 22701 814 22735
rect 848 22701 877 22735
rect 757 22663 877 22701
rect 757 22629 814 22663
rect 848 22629 877 22663
rect 757 22591 877 22629
rect 757 22557 814 22591
rect 848 22557 877 22591
rect 757 22519 877 22557
rect 757 22485 814 22519
rect 848 22485 877 22519
rect 757 22447 877 22485
rect 757 22413 814 22447
rect 848 22413 877 22447
rect 757 22375 877 22413
rect 757 22341 814 22375
rect 848 22341 877 22375
rect 757 22303 877 22341
rect 757 22269 814 22303
rect 848 22269 877 22303
rect 757 22231 877 22269
rect 757 22197 814 22231
rect 848 22197 877 22231
rect 757 22159 877 22197
rect 757 22125 814 22159
rect 848 22125 877 22159
rect 757 22087 877 22125
rect 757 22053 814 22087
rect 848 22053 877 22087
rect 757 22015 877 22053
rect 757 21981 814 22015
rect 848 21981 877 22015
rect 757 21943 877 21981
rect 757 21909 814 21943
rect 848 21909 877 21943
rect 757 21871 877 21909
rect 757 21837 814 21871
rect 848 21837 877 21871
rect 757 21799 877 21837
rect 757 21765 814 21799
rect 848 21765 877 21799
rect 757 21727 877 21765
rect 757 21693 814 21727
rect 848 21693 877 21727
rect 757 21655 877 21693
rect 757 21621 814 21655
rect 848 21621 877 21655
rect 757 21583 877 21621
rect 757 21549 814 21583
rect 848 21549 877 21583
rect 757 21511 877 21549
rect 757 21477 814 21511
rect 848 21477 877 21511
rect 757 21439 877 21477
rect 757 21405 814 21439
rect 848 21405 877 21439
rect 757 21367 877 21405
rect 757 21333 814 21367
rect 848 21333 877 21367
rect 757 21295 877 21333
rect 757 21261 814 21295
rect 848 21261 877 21295
rect 757 21223 877 21261
rect 757 21189 814 21223
rect 848 21189 877 21223
rect 757 21151 877 21189
rect 757 21117 814 21151
rect 848 21117 877 21151
rect 757 21079 877 21117
rect 757 21045 814 21079
rect 848 21045 877 21079
rect 757 21007 877 21045
rect 757 20973 814 21007
rect 848 20973 877 21007
rect 757 20935 877 20973
rect 757 20901 814 20935
rect 848 20901 877 20935
rect 757 20863 877 20901
rect 757 20829 814 20863
rect 848 20829 877 20863
rect 757 20791 877 20829
rect 757 20757 814 20791
rect 848 20757 877 20791
rect 757 20719 877 20757
rect 757 20685 814 20719
rect 848 20685 877 20719
rect 757 20647 877 20685
rect 757 20613 814 20647
rect 848 20613 877 20647
rect 757 20575 877 20613
rect 757 20541 814 20575
rect 848 20541 877 20575
rect 757 20503 877 20541
rect 757 20469 814 20503
rect 848 20469 877 20503
rect 757 20431 877 20469
rect 757 20397 814 20431
rect 848 20397 877 20431
rect 757 20359 877 20397
rect 757 20325 814 20359
rect 848 20325 877 20359
rect 757 20287 877 20325
rect 757 20253 814 20287
rect 848 20253 877 20287
rect 757 20215 877 20253
rect 757 20181 814 20215
rect 848 20181 877 20215
rect 757 20143 877 20181
rect 757 20109 814 20143
rect 848 20109 877 20143
rect 757 20071 877 20109
rect 757 20037 814 20071
rect 848 20037 877 20071
rect 757 19999 877 20037
rect 757 19965 814 19999
rect 848 19965 877 19999
rect 757 19927 877 19965
rect 757 19893 814 19927
rect 848 19893 877 19927
rect 757 19855 877 19893
rect 757 19821 814 19855
rect 848 19821 877 19855
rect 757 19783 877 19821
rect 757 19749 814 19783
rect 848 19749 877 19783
rect 757 19711 877 19749
rect 757 19677 814 19711
rect 848 19677 877 19711
rect 757 19639 877 19677
rect 757 19605 814 19639
rect 848 19605 877 19639
rect 757 19567 877 19605
rect 757 19533 814 19567
rect 848 19533 877 19567
rect 757 19495 877 19533
rect 757 19461 814 19495
rect 848 19461 877 19495
rect 757 19423 877 19461
rect 757 19389 814 19423
rect 848 19389 877 19423
rect 757 19351 877 19389
rect 757 19317 814 19351
rect 848 19317 877 19351
rect 757 19279 877 19317
rect 757 19245 814 19279
rect 848 19245 877 19279
rect 757 19207 877 19245
rect 757 19173 814 19207
rect 848 19173 877 19207
rect 757 19135 877 19173
rect 757 19101 814 19135
rect 848 19101 877 19135
rect 757 19063 877 19101
rect 757 19029 814 19063
rect 848 19029 877 19063
rect 757 18991 877 19029
rect 757 18957 814 18991
rect 848 18957 877 18991
rect 757 18919 877 18957
rect 757 18885 814 18919
rect 848 18885 877 18919
rect 757 18847 877 18885
rect 757 18813 814 18847
rect 848 18813 877 18847
rect 757 18775 877 18813
rect 757 18741 814 18775
rect 848 18741 877 18775
rect 757 18703 877 18741
rect 757 18669 814 18703
rect 848 18669 877 18703
rect 757 18631 877 18669
rect 757 18597 814 18631
rect 848 18597 877 18631
rect 757 18559 877 18597
rect 757 18525 814 18559
rect 848 18525 877 18559
rect 757 18487 877 18525
rect 757 18453 814 18487
rect 848 18453 877 18487
rect 757 18415 877 18453
rect 757 18381 814 18415
rect 848 18381 877 18415
rect 757 18343 877 18381
rect 757 18309 814 18343
rect 848 18309 877 18343
rect 757 18271 877 18309
rect 757 18237 814 18271
rect 848 18237 877 18271
rect 757 18199 877 18237
rect 757 18165 814 18199
rect 848 18165 877 18199
rect 757 18127 877 18165
rect 757 18093 814 18127
rect 848 18093 877 18127
rect 757 18055 877 18093
rect 757 18021 814 18055
rect 848 18021 877 18055
rect 757 17983 877 18021
rect 757 17949 814 17983
rect 848 17949 877 17983
rect 757 17911 877 17949
rect 757 17877 814 17911
rect 848 17877 877 17911
rect 757 17839 877 17877
rect 757 17805 814 17839
rect 848 17805 877 17839
rect 757 17767 877 17805
rect 757 17733 814 17767
rect 848 17733 877 17767
rect 757 17695 877 17733
rect 757 17661 814 17695
rect 848 17661 877 17695
rect 757 17623 877 17661
rect 757 17589 814 17623
rect 848 17589 877 17623
rect 757 17551 877 17589
rect 757 17517 814 17551
rect 848 17517 877 17551
rect 757 17479 877 17517
rect 757 17445 814 17479
rect 848 17445 877 17479
rect 757 17407 877 17445
rect 757 17373 814 17407
rect 848 17373 877 17407
rect 757 17335 877 17373
rect 757 17301 814 17335
rect 848 17301 877 17335
rect 757 17263 877 17301
rect 757 17229 814 17263
rect 848 17229 877 17263
rect 757 17191 877 17229
rect 757 17157 814 17191
rect 848 17157 877 17191
rect 757 17119 877 17157
rect 757 17085 814 17119
rect 848 17085 877 17119
rect 757 17047 877 17085
rect 757 17013 814 17047
rect 848 17013 877 17047
rect 757 16975 877 17013
rect 757 16941 814 16975
rect 848 16941 877 16975
rect 757 16903 877 16941
rect 757 16869 814 16903
rect 848 16869 877 16903
rect 757 16831 877 16869
rect 757 16797 814 16831
rect 848 16797 877 16831
rect 757 16759 877 16797
rect 757 16725 814 16759
rect 848 16725 877 16759
rect 757 16687 877 16725
rect 757 16653 814 16687
rect 848 16653 877 16687
rect 757 16615 877 16653
rect 757 16581 814 16615
rect 848 16581 877 16615
rect 757 16543 877 16581
rect 757 16509 814 16543
rect 848 16509 877 16543
rect 757 16471 877 16509
rect 757 16437 814 16471
rect 848 16437 877 16471
rect 757 16399 877 16437
rect 757 16365 814 16399
rect 848 16365 877 16399
rect 757 16327 877 16365
rect 757 16293 814 16327
rect 848 16293 877 16327
rect 757 16255 877 16293
rect 757 16221 814 16255
rect 848 16221 877 16255
rect 757 16183 877 16221
rect 757 16149 814 16183
rect 848 16149 877 16183
rect 757 16111 877 16149
rect 757 16077 814 16111
rect 848 16077 877 16111
rect 757 16039 877 16077
rect 757 16005 814 16039
rect 848 16005 877 16039
rect 757 15967 877 16005
rect 757 15933 814 15967
rect 848 15933 877 15967
rect 757 15895 877 15933
rect 757 15861 814 15895
rect 848 15861 877 15895
rect 757 15823 877 15861
rect 757 15789 814 15823
rect 848 15789 877 15823
rect 757 15751 877 15789
rect 757 15717 814 15751
rect 848 15717 877 15751
rect 757 15679 877 15717
rect 757 15645 814 15679
rect 848 15645 877 15679
rect 757 15607 877 15645
rect 757 15573 814 15607
rect 848 15573 877 15607
rect 757 15535 877 15573
rect 757 15501 814 15535
rect 848 15501 877 15535
rect 757 15463 877 15501
rect 757 15429 814 15463
rect 848 15429 877 15463
rect 757 15391 877 15429
rect 757 15357 814 15391
rect 848 15357 877 15391
rect 757 15319 877 15357
rect 757 15285 814 15319
rect 848 15285 877 15319
rect 757 15247 877 15285
rect 757 15213 814 15247
rect 848 15213 877 15247
rect 757 15175 877 15213
rect 757 15141 814 15175
rect 848 15141 877 15175
rect 757 15103 877 15141
rect 757 15069 814 15103
rect 848 15069 877 15103
rect 757 15031 877 15069
rect 757 14997 814 15031
rect 848 14997 877 15031
rect 757 14959 877 14997
rect 757 14925 814 14959
rect 848 14925 877 14959
rect 757 14887 877 14925
rect 757 14853 814 14887
rect 848 14853 877 14887
rect 757 14815 877 14853
rect 757 14781 814 14815
rect 848 14781 877 14815
rect 757 14743 877 14781
rect 757 14709 814 14743
rect 848 14709 877 14743
rect 757 14671 877 14709
rect 757 14637 814 14671
rect 848 14637 877 14671
rect 757 14599 877 14637
rect 757 14565 814 14599
rect 848 14565 877 14599
rect 757 14527 877 14565
rect 757 14493 814 14527
rect 848 14493 877 14527
rect 757 14455 877 14493
rect 757 14421 814 14455
rect 848 14421 877 14455
rect 757 14383 877 14421
rect 757 14349 814 14383
rect 848 14349 877 14383
rect 757 14311 877 14349
rect 757 14277 814 14311
rect 848 14277 877 14311
rect 757 14239 877 14277
rect 757 14205 814 14239
rect 848 14205 877 14239
rect 757 14167 877 14205
rect 757 14133 814 14167
rect 848 14133 877 14167
rect 757 14095 877 14133
rect 757 14061 814 14095
rect 848 14061 877 14095
rect 757 14023 877 14061
rect 757 13989 814 14023
rect 848 13989 877 14023
rect 757 13951 877 13989
rect 757 13917 814 13951
rect 848 13917 877 13951
rect 757 13879 877 13917
rect 757 13845 814 13879
rect 848 13845 877 13879
rect 757 13807 877 13845
rect 757 13773 814 13807
rect 848 13773 877 13807
rect 757 13735 877 13773
rect 757 13701 814 13735
rect 848 13701 877 13735
rect 757 13663 877 13701
rect 757 13629 814 13663
rect 848 13629 877 13663
rect 757 13591 877 13629
rect 757 13557 814 13591
rect 848 13557 877 13591
rect 757 13519 877 13557
rect 757 13485 814 13519
rect 848 13485 877 13519
rect 757 13447 877 13485
rect 757 13413 814 13447
rect 848 13413 877 13447
rect 757 13375 877 13413
rect 757 13341 814 13375
rect 848 13341 877 13375
rect 757 13303 877 13341
rect 757 13269 814 13303
rect 848 13269 877 13303
rect 757 13231 877 13269
rect 757 13197 814 13231
rect 848 13197 877 13231
rect 757 13159 877 13197
rect 757 13125 814 13159
rect 848 13125 877 13159
rect 757 13087 877 13125
rect 757 13053 814 13087
rect 848 13053 877 13087
rect 757 13015 877 13053
rect 757 12981 814 13015
rect 848 12981 877 13015
rect 757 12943 877 12981
rect 757 12909 814 12943
rect 848 12909 877 12943
rect 757 12871 877 12909
rect 757 12837 814 12871
rect 848 12837 877 12871
rect 757 12799 877 12837
rect 757 12765 814 12799
rect 848 12765 877 12799
rect 757 12727 877 12765
rect 757 12693 814 12727
rect 848 12693 877 12727
rect 757 12655 877 12693
rect 757 12621 814 12655
rect 848 12621 877 12655
rect 757 12583 877 12621
rect 757 12549 814 12583
rect 848 12549 877 12583
rect 757 12511 877 12549
rect 757 12477 814 12511
rect 848 12477 877 12511
rect 757 12439 877 12477
rect 757 12405 814 12439
rect 848 12405 877 12439
rect 757 12367 877 12405
rect 757 12333 814 12367
rect 848 12333 877 12367
rect 757 12295 877 12333
rect 757 12261 814 12295
rect 848 12261 877 12295
rect 757 12223 877 12261
rect 757 12189 814 12223
rect 848 12189 877 12223
rect 757 12151 877 12189
rect 757 12117 814 12151
rect 848 12117 877 12151
rect 757 12079 877 12117
rect 757 12045 814 12079
rect 848 12045 877 12079
rect 757 12007 877 12045
rect 757 11973 814 12007
rect 848 11973 877 12007
rect 757 11935 877 11973
rect 757 11901 814 11935
rect 848 11901 877 11935
rect 757 11863 877 11901
rect 757 11829 814 11863
rect 848 11829 877 11863
rect 757 11791 877 11829
rect 757 11757 814 11791
rect 848 11757 877 11791
rect 757 11719 877 11757
rect 757 11685 814 11719
rect 848 11685 877 11719
rect 757 11647 877 11685
rect 757 11613 814 11647
rect 848 11613 877 11647
rect 757 11575 877 11613
rect 757 11541 814 11575
rect 848 11541 877 11575
rect 757 11503 877 11541
rect 757 11469 814 11503
rect 848 11469 877 11503
rect 757 11431 877 11469
rect 757 11397 814 11431
rect 848 11397 877 11431
rect 757 11359 877 11397
rect 757 11325 814 11359
rect 848 11325 877 11359
rect 757 11287 877 11325
rect 757 11253 814 11287
rect 848 11253 877 11287
rect 757 11215 877 11253
rect 757 11181 814 11215
rect 848 11181 877 11215
rect 757 11143 877 11181
rect 757 11109 814 11143
rect 848 11109 877 11143
rect 757 11071 877 11109
rect 757 11037 814 11071
rect 848 11037 877 11071
rect 757 10999 877 11037
rect 757 10965 814 10999
rect 848 10965 877 10999
rect 757 10927 877 10965
rect 757 10893 814 10927
rect 848 10893 877 10927
rect 757 10855 877 10893
rect 757 10821 814 10855
rect 848 10821 877 10855
rect 757 10783 877 10821
rect 757 10749 814 10783
rect 848 10749 877 10783
rect 757 10711 877 10749
rect 757 10677 814 10711
rect 848 10677 877 10711
rect 757 10639 877 10677
rect 757 10605 814 10639
rect 848 10605 877 10639
rect 757 10567 877 10605
rect 757 10533 814 10567
rect 848 10533 877 10567
rect 757 10495 877 10533
rect 757 10461 814 10495
rect 848 10461 877 10495
rect 757 10423 877 10461
rect 757 10389 814 10423
rect 848 10389 877 10423
rect 757 10351 877 10389
rect 757 10317 814 10351
rect 848 10317 877 10351
rect 757 10279 877 10317
rect 757 10245 814 10279
rect 848 10245 877 10279
rect 757 10207 877 10245
rect 1177 34636 13817 34684
rect 1177 34602 1365 34636
rect 1399 34602 1437 34636
rect 1471 34602 1509 34636
rect 1543 34602 1581 34636
rect 1615 34602 1653 34636
rect 1687 34602 1725 34636
rect 1759 34602 1797 34636
rect 1831 34602 1869 34636
rect 1903 34602 1941 34636
rect 1975 34602 2013 34636
rect 2047 34602 2085 34636
rect 2119 34602 2157 34636
rect 2191 34602 2229 34636
rect 2263 34602 2301 34636
rect 2335 34602 2373 34636
rect 2407 34602 2445 34636
rect 2479 34602 2517 34636
rect 2551 34602 2589 34636
rect 2623 34602 2661 34636
rect 2695 34602 2733 34636
rect 2767 34602 2805 34636
rect 2839 34602 2877 34636
rect 2911 34602 2949 34636
rect 2983 34602 3021 34636
rect 3055 34602 3093 34636
rect 3127 34602 3165 34636
rect 3199 34602 3237 34636
rect 3271 34602 3309 34636
rect 3343 34602 3381 34636
rect 3415 34602 3453 34636
rect 3487 34602 3525 34636
rect 3559 34602 3597 34636
rect 3631 34602 3669 34636
rect 3703 34602 3741 34636
rect 3775 34602 3813 34636
rect 3847 34602 3885 34636
rect 3919 34602 3957 34636
rect 3991 34602 4029 34636
rect 4063 34602 4101 34636
rect 4135 34602 4173 34636
rect 4207 34602 4245 34636
rect 4279 34602 4317 34636
rect 4351 34602 4389 34636
rect 4423 34602 4461 34636
rect 4495 34602 4533 34636
rect 4567 34602 4605 34636
rect 4639 34602 4677 34636
rect 4711 34602 4749 34636
rect 4783 34602 4821 34636
rect 4855 34602 4893 34636
rect 4927 34602 4965 34636
rect 4999 34602 5037 34636
rect 5071 34602 5109 34636
rect 5143 34602 5181 34636
rect 5215 34602 5253 34636
rect 5287 34602 5325 34636
rect 5359 34602 5397 34636
rect 5431 34602 5469 34636
rect 5503 34602 5541 34636
rect 5575 34602 5613 34636
rect 5647 34602 5685 34636
rect 5719 34602 5757 34636
rect 5791 34602 5829 34636
rect 5863 34602 5901 34636
rect 5935 34602 5973 34636
rect 6007 34602 6045 34636
rect 6079 34602 6117 34636
rect 6151 34602 6189 34636
rect 6223 34602 6261 34636
rect 6295 34602 6333 34636
rect 6367 34602 6405 34636
rect 6439 34602 6477 34636
rect 6511 34602 6549 34636
rect 6583 34602 6621 34636
rect 6655 34602 6693 34636
rect 6727 34602 6765 34636
rect 6799 34602 6837 34636
rect 6871 34602 6909 34636
rect 6943 34602 6981 34636
rect 7015 34602 7053 34636
rect 7087 34602 7125 34636
rect 7159 34602 7197 34636
rect 7231 34602 7269 34636
rect 7303 34602 7341 34636
rect 7375 34602 7413 34636
rect 7447 34602 7485 34636
rect 7519 34602 7557 34636
rect 7591 34602 7629 34636
rect 7663 34602 7701 34636
rect 7735 34602 7773 34636
rect 7807 34602 7845 34636
rect 7879 34602 7917 34636
rect 7951 34602 7989 34636
rect 8023 34602 8061 34636
rect 8095 34602 8133 34636
rect 8167 34602 8205 34636
rect 8239 34602 8277 34636
rect 8311 34602 8349 34636
rect 8383 34602 8421 34636
rect 8455 34602 8493 34636
rect 8527 34602 8565 34636
rect 8599 34602 8637 34636
rect 8671 34602 8709 34636
rect 8743 34602 8781 34636
rect 8815 34602 8853 34636
rect 8887 34602 8925 34636
rect 8959 34602 8997 34636
rect 9031 34602 9069 34636
rect 9103 34602 9141 34636
rect 9175 34602 9213 34636
rect 9247 34602 9285 34636
rect 9319 34602 9357 34636
rect 9391 34602 9429 34636
rect 9463 34602 9501 34636
rect 9535 34602 9573 34636
rect 9607 34602 9645 34636
rect 9679 34602 9717 34636
rect 9751 34602 9789 34636
rect 9823 34602 9861 34636
rect 9895 34602 9933 34636
rect 9967 34602 10005 34636
rect 10039 34602 10077 34636
rect 10111 34602 10149 34636
rect 10183 34602 10221 34636
rect 10255 34602 10293 34636
rect 10327 34602 10365 34636
rect 10399 34602 10437 34636
rect 10471 34602 10509 34636
rect 10543 34602 10581 34636
rect 10615 34602 10653 34636
rect 10687 34602 10725 34636
rect 10759 34602 10797 34636
rect 10831 34602 10869 34636
rect 10903 34602 10941 34636
rect 10975 34602 11013 34636
rect 11047 34602 11085 34636
rect 11119 34602 11157 34636
rect 11191 34602 11229 34636
rect 11263 34602 11301 34636
rect 11335 34602 11373 34636
rect 11407 34602 11445 34636
rect 11479 34602 11517 34636
rect 11551 34602 11589 34636
rect 11623 34602 11661 34636
rect 11695 34602 11733 34636
rect 11767 34602 11805 34636
rect 11839 34602 11877 34636
rect 11911 34602 11949 34636
rect 11983 34602 12021 34636
rect 12055 34602 12093 34636
rect 12127 34602 12165 34636
rect 12199 34602 12237 34636
rect 12271 34602 12309 34636
rect 12343 34602 12381 34636
rect 12415 34602 12453 34636
rect 12487 34602 12525 34636
rect 12559 34602 12597 34636
rect 12631 34602 12669 34636
rect 12703 34602 12741 34636
rect 12775 34602 12813 34636
rect 12847 34602 12885 34636
rect 12919 34602 12957 34636
rect 12991 34602 13029 34636
rect 13063 34602 13101 34636
rect 13135 34602 13173 34636
rect 13207 34602 13245 34636
rect 13279 34602 13317 34636
rect 13351 34602 13389 34636
rect 13423 34602 13461 34636
rect 13495 34602 13533 34636
rect 13567 34602 13605 34636
rect 13639 34602 13817 34636
rect 1177 34564 13817 34602
rect 1177 34474 1297 34564
rect 1177 34440 1221 34474
rect 1255 34440 1297 34474
rect 1177 34402 1297 34440
rect 1177 34368 1221 34402
rect 1255 34368 1297 34402
rect 1177 34330 1297 34368
rect 1177 34296 1221 34330
rect 1255 34296 1297 34330
rect 1177 34258 1297 34296
rect 1177 34224 1221 34258
rect 1255 34224 1297 34258
rect 1177 34186 1297 34224
rect 1177 34152 1221 34186
rect 1255 34152 1297 34186
rect 1177 34114 1297 34152
rect 1177 34080 1221 34114
rect 1255 34080 1297 34114
rect 1177 34042 1297 34080
rect 1177 34008 1221 34042
rect 1255 34008 1297 34042
rect 1177 33970 1297 34008
rect 1177 33936 1221 33970
rect 1255 33936 1297 33970
rect 1177 33898 1297 33936
rect 1177 33864 1221 33898
rect 1255 33864 1297 33898
rect 1177 33826 1297 33864
rect 1177 33792 1221 33826
rect 1255 33792 1297 33826
rect 1177 33754 1297 33792
rect 1177 33720 1221 33754
rect 1255 33720 1297 33754
rect 1177 33682 1297 33720
rect 1177 33648 1221 33682
rect 1255 33648 1297 33682
rect 1177 33610 1297 33648
rect 1177 33576 1221 33610
rect 1255 33576 1297 33610
rect 1177 33538 1297 33576
rect 1177 33504 1221 33538
rect 1255 33504 1297 33538
rect 1177 33466 1297 33504
rect 1177 33432 1221 33466
rect 1255 33432 1297 33466
rect 1177 33394 1297 33432
rect 1177 33360 1221 33394
rect 1255 33360 1297 33394
rect 1177 33322 1297 33360
rect 1177 33288 1221 33322
rect 1255 33288 1297 33322
rect 1177 33250 1297 33288
rect 1177 33216 1221 33250
rect 1255 33216 1297 33250
rect 1177 33178 1297 33216
rect 1177 33144 1221 33178
rect 1255 33144 1297 33178
rect 1177 33106 1297 33144
rect 1177 33072 1221 33106
rect 1255 33072 1297 33106
rect 1177 33034 1297 33072
rect 1177 33000 1221 33034
rect 1255 33000 1297 33034
rect 1177 32962 1297 33000
rect 1177 32928 1221 32962
rect 1255 32928 1297 32962
rect 1177 32890 1297 32928
rect 1177 32856 1221 32890
rect 1255 32856 1297 32890
rect 1177 32818 1297 32856
rect 1177 32784 1221 32818
rect 1255 32784 1297 32818
rect 1177 32746 1297 32784
rect 1177 32712 1221 32746
rect 1255 32712 1297 32746
rect 1177 32674 1297 32712
rect 1177 32640 1221 32674
rect 1255 32640 1297 32674
rect 1177 32602 1297 32640
rect 1177 32568 1221 32602
rect 1255 32568 1297 32602
rect 1177 32530 1297 32568
rect 1177 32496 1221 32530
rect 1255 32496 1297 32530
rect 1177 32458 1297 32496
rect 1177 32424 1221 32458
rect 1255 32424 1297 32458
rect 1177 32386 1297 32424
rect 1177 32352 1221 32386
rect 1255 32352 1297 32386
rect 1177 32314 1297 32352
rect 1177 32280 1221 32314
rect 1255 32280 1297 32314
rect 1177 32242 1297 32280
rect 1177 32208 1221 32242
rect 1255 32208 1297 32242
rect 1177 32170 1297 32208
rect 1177 32136 1221 32170
rect 1255 32136 1297 32170
rect 1177 32098 1297 32136
rect 1177 32064 1221 32098
rect 1255 32064 1297 32098
rect 1177 32026 1297 32064
rect 1177 31992 1221 32026
rect 1255 31992 1297 32026
rect 1177 31954 1297 31992
rect 1177 31920 1221 31954
rect 1255 31920 1297 31954
rect 1177 31882 1297 31920
rect 1177 31848 1221 31882
rect 1255 31848 1297 31882
rect 1177 31810 1297 31848
rect 1177 31776 1221 31810
rect 1255 31776 1297 31810
rect 1177 31738 1297 31776
rect 1177 31704 1221 31738
rect 1255 31704 1297 31738
rect 1177 31666 1297 31704
rect 1177 31632 1221 31666
rect 1255 31632 1297 31666
rect 1177 31594 1297 31632
rect 1177 31560 1221 31594
rect 1255 31560 1297 31594
rect 1177 31522 1297 31560
rect 1177 31488 1221 31522
rect 1255 31488 1297 31522
rect 1177 31450 1297 31488
rect 1177 31416 1221 31450
rect 1255 31416 1297 31450
rect 1177 31378 1297 31416
rect 1177 31344 1221 31378
rect 1255 31344 1297 31378
rect 1177 31306 1297 31344
rect 1177 31272 1221 31306
rect 1255 31272 1297 31306
rect 1177 31234 1297 31272
rect 1177 31200 1221 31234
rect 1255 31200 1297 31234
rect 1177 31162 1297 31200
rect 1177 31128 1221 31162
rect 1255 31128 1297 31162
rect 1177 31090 1297 31128
rect 1177 31056 1221 31090
rect 1255 31056 1297 31090
rect 1177 31018 1297 31056
rect 1177 30984 1221 31018
rect 1255 30984 1297 31018
rect 1177 30946 1297 30984
rect 1177 30912 1221 30946
rect 1255 30912 1297 30946
rect 1177 30874 1297 30912
rect 1177 30840 1221 30874
rect 1255 30840 1297 30874
rect 1177 30802 1297 30840
rect 1177 30768 1221 30802
rect 1255 30768 1297 30802
rect 1177 30730 1297 30768
rect 1177 30696 1221 30730
rect 1255 30696 1297 30730
rect 1177 30658 1297 30696
rect 1177 30624 1221 30658
rect 1255 30624 1297 30658
rect 1177 30586 1297 30624
rect 1177 30552 1221 30586
rect 1255 30552 1297 30586
rect 1177 30514 1297 30552
rect 1177 30480 1221 30514
rect 1255 30480 1297 30514
rect 1177 30442 1297 30480
rect 1177 30408 1221 30442
rect 1255 30408 1297 30442
rect 1177 30370 1297 30408
rect 1177 30336 1221 30370
rect 1255 30336 1297 30370
rect 1177 30298 1297 30336
rect 1177 30264 1221 30298
rect 1255 30264 1297 30298
rect 1177 30226 1297 30264
rect 1177 30192 1221 30226
rect 1255 30192 1297 30226
rect 1177 30154 1297 30192
rect 1177 30120 1221 30154
rect 1255 30120 1297 30154
rect 1177 30082 1297 30120
rect 1177 30048 1221 30082
rect 1255 30048 1297 30082
rect 1177 30010 1297 30048
rect 1177 29976 1221 30010
rect 1255 29976 1297 30010
rect 1177 29938 1297 29976
rect 1177 29904 1221 29938
rect 1255 29904 1297 29938
rect 1177 29866 1297 29904
rect 1177 29832 1221 29866
rect 1255 29832 1297 29866
rect 1177 29794 1297 29832
rect 1177 29760 1221 29794
rect 1255 29760 1297 29794
rect 1177 29722 1297 29760
rect 1177 29688 1221 29722
rect 1255 29688 1297 29722
rect 1177 29650 1297 29688
rect 1177 29616 1221 29650
rect 1255 29616 1297 29650
rect 1177 29578 1297 29616
rect 1177 29544 1221 29578
rect 1255 29544 1297 29578
rect 1177 29506 1297 29544
rect 1177 29472 1221 29506
rect 1255 29472 1297 29506
rect 1177 29434 1297 29472
rect 1177 29400 1221 29434
rect 1255 29400 1297 29434
rect 1177 29362 1297 29400
rect 1177 29328 1221 29362
rect 1255 29328 1297 29362
rect 1177 29290 1297 29328
rect 1177 29256 1221 29290
rect 1255 29256 1297 29290
rect 1177 29218 1297 29256
rect 1177 29184 1221 29218
rect 1255 29184 1297 29218
rect 1177 29146 1297 29184
rect 1177 29112 1221 29146
rect 1255 29112 1297 29146
rect 1177 29074 1297 29112
rect 1177 29040 1221 29074
rect 1255 29040 1297 29074
rect 1177 29002 1297 29040
rect 1177 28968 1221 29002
rect 1255 28968 1297 29002
rect 1177 28930 1297 28968
rect 1177 28896 1221 28930
rect 1255 28896 1297 28930
rect 1177 28858 1297 28896
rect 1177 28824 1221 28858
rect 1255 28824 1297 28858
rect 1177 28786 1297 28824
rect 1177 28752 1221 28786
rect 1255 28752 1297 28786
rect 1177 28714 1297 28752
rect 1177 28680 1221 28714
rect 1255 28680 1297 28714
rect 1177 28642 1297 28680
rect 1177 28608 1221 28642
rect 1255 28608 1297 28642
rect 1177 28570 1297 28608
rect 1177 28536 1221 28570
rect 1255 28536 1297 28570
rect 1177 28498 1297 28536
rect 1177 28464 1221 28498
rect 1255 28464 1297 28498
rect 1177 28426 1297 28464
rect 1177 28392 1221 28426
rect 1255 28392 1297 28426
rect 1177 28354 1297 28392
rect 1177 28320 1221 28354
rect 1255 28320 1297 28354
rect 1177 28282 1297 28320
rect 1177 28248 1221 28282
rect 1255 28248 1297 28282
rect 1177 28210 1297 28248
rect 1177 28176 1221 28210
rect 1255 28176 1297 28210
rect 1177 28138 1297 28176
rect 1177 28104 1221 28138
rect 1255 28104 1297 28138
rect 1177 28066 1297 28104
rect 1177 28032 1221 28066
rect 1255 28032 1297 28066
rect 1177 27994 1297 28032
rect 1177 27960 1221 27994
rect 1255 27960 1297 27994
rect 1177 27922 1297 27960
rect 1177 27888 1221 27922
rect 1255 27888 1297 27922
rect 1177 27850 1297 27888
rect 1177 27816 1221 27850
rect 1255 27816 1297 27850
rect 1177 27778 1297 27816
rect 1177 27744 1221 27778
rect 1255 27744 1297 27778
rect 1177 27706 1297 27744
rect 1177 27672 1221 27706
rect 1255 27672 1297 27706
rect 1177 27634 1297 27672
rect 1177 27600 1221 27634
rect 1255 27600 1297 27634
rect 1177 27562 1297 27600
rect 1177 27528 1221 27562
rect 1255 27528 1297 27562
rect 1177 27490 1297 27528
rect 1177 27456 1221 27490
rect 1255 27456 1297 27490
rect 1177 27418 1297 27456
rect 1177 27384 1221 27418
rect 1255 27384 1297 27418
rect 1177 27346 1297 27384
rect 1177 27312 1221 27346
rect 1255 27312 1297 27346
rect 1177 27274 1297 27312
rect 1177 27240 1221 27274
rect 1255 27240 1297 27274
rect 1177 27202 1297 27240
rect 1177 27168 1221 27202
rect 1255 27168 1297 27202
rect 1177 27130 1297 27168
rect 1177 27096 1221 27130
rect 1255 27096 1297 27130
rect 1177 27058 1297 27096
rect 1177 27024 1221 27058
rect 1255 27024 1297 27058
rect 1177 26986 1297 27024
rect 1177 26952 1221 26986
rect 1255 26952 1297 26986
rect 1177 26914 1297 26952
rect 1177 26880 1221 26914
rect 1255 26880 1297 26914
rect 1177 26842 1297 26880
rect 1177 26808 1221 26842
rect 1255 26808 1297 26842
rect 1177 26770 1297 26808
rect 1177 26736 1221 26770
rect 1255 26736 1297 26770
rect 1177 26698 1297 26736
rect 1177 26664 1221 26698
rect 1255 26664 1297 26698
rect 1177 26626 1297 26664
rect 1177 26592 1221 26626
rect 1255 26592 1297 26626
rect 1177 26554 1297 26592
rect 1177 26520 1221 26554
rect 1255 26520 1297 26554
rect 1177 26482 1297 26520
rect 1177 26448 1221 26482
rect 1255 26448 1297 26482
rect 1177 26410 1297 26448
rect 1177 26376 1221 26410
rect 1255 26376 1297 26410
rect 1177 26338 1297 26376
rect 1177 26304 1221 26338
rect 1255 26304 1297 26338
rect 1177 26266 1297 26304
rect 1177 26232 1221 26266
rect 1255 26232 1297 26266
rect 1177 26194 1297 26232
rect 1177 26160 1221 26194
rect 1255 26160 1297 26194
rect 1177 26122 1297 26160
rect 1177 26088 1221 26122
rect 1255 26088 1297 26122
rect 1177 26050 1297 26088
rect 1177 26016 1221 26050
rect 1255 26016 1297 26050
rect 1177 25978 1297 26016
rect 1177 25944 1221 25978
rect 1255 25944 1297 25978
rect 1177 25906 1297 25944
rect 1177 25872 1221 25906
rect 1255 25872 1297 25906
rect 1177 25834 1297 25872
rect 1177 25800 1221 25834
rect 1255 25800 1297 25834
rect 1177 25762 1297 25800
rect 1177 25728 1221 25762
rect 1255 25728 1297 25762
rect 1177 25690 1297 25728
rect 1177 25656 1221 25690
rect 1255 25656 1297 25690
rect 1177 25618 1297 25656
rect 1177 25584 1221 25618
rect 1255 25584 1297 25618
rect 1177 25546 1297 25584
rect 1177 25512 1221 25546
rect 1255 25512 1297 25546
rect 1177 25474 1297 25512
rect 1177 25440 1221 25474
rect 1255 25440 1297 25474
rect 1177 25402 1297 25440
rect 1177 25368 1221 25402
rect 1255 25368 1297 25402
rect 1177 25330 1297 25368
rect 1177 25296 1221 25330
rect 1255 25296 1297 25330
rect 1177 25258 1297 25296
rect 1177 25224 1221 25258
rect 1255 25224 1297 25258
rect 1177 25186 1297 25224
rect 1177 25152 1221 25186
rect 1255 25152 1297 25186
rect 1177 25114 1297 25152
rect 1177 25080 1221 25114
rect 1255 25080 1297 25114
rect 1177 25042 1297 25080
rect 1177 25008 1221 25042
rect 1255 25008 1297 25042
rect 1177 24970 1297 25008
rect 1177 24936 1221 24970
rect 1255 24936 1297 24970
rect 1177 24898 1297 24936
rect 1177 24864 1221 24898
rect 1255 24864 1297 24898
rect 1177 24826 1297 24864
rect 1177 24792 1221 24826
rect 1255 24792 1297 24826
rect 1177 24754 1297 24792
rect 1177 24720 1221 24754
rect 1255 24720 1297 24754
rect 1177 24682 1297 24720
rect 1177 24648 1221 24682
rect 1255 24648 1297 24682
rect 1177 24610 1297 24648
rect 1177 24576 1221 24610
rect 1255 24576 1297 24610
rect 1177 24538 1297 24576
rect 1177 24504 1221 24538
rect 1255 24504 1297 24538
rect 1177 24466 1297 24504
rect 1177 24432 1221 24466
rect 1255 24432 1297 24466
rect 1177 24394 1297 24432
rect 1177 24360 1221 24394
rect 1255 24360 1297 24394
rect 1177 24322 1297 24360
rect 1177 24288 1221 24322
rect 1255 24288 1297 24322
rect 1177 24250 1297 24288
rect 1177 24216 1221 24250
rect 1255 24216 1297 24250
rect 1177 24178 1297 24216
rect 1177 24144 1221 24178
rect 1255 24144 1297 24178
rect 1177 24106 1297 24144
rect 1177 24072 1221 24106
rect 1255 24072 1297 24106
rect 1177 24034 1297 24072
rect 1177 24000 1221 24034
rect 1255 24000 1297 24034
rect 1177 23962 1297 24000
rect 1177 23928 1221 23962
rect 1255 23928 1297 23962
rect 1177 23890 1297 23928
rect 1177 23856 1221 23890
rect 1255 23856 1297 23890
rect 1177 23818 1297 23856
rect 1177 23784 1221 23818
rect 1255 23784 1297 23818
rect 1177 23746 1297 23784
rect 1177 23712 1221 23746
rect 1255 23712 1297 23746
rect 1177 23674 1297 23712
rect 1177 23640 1221 23674
rect 1255 23640 1297 23674
rect 1177 23602 1297 23640
rect 1177 23568 1221 23602
rect 1255 23568 1297 23602
rect 1177 23530 1297 23568
rect 1177 23496 1221 23530
rect 1255 23496 1297 23530
rect 1177 23458 1297 23496
rect 1177 23424 1221 23458
rect 1255 23424 1297 23458
rect 1177 23386 1297 23424
rect 1177 23352 1221 23386
rect 1255 23352 1297 23386
rect 1177 23314 1297 23352
rect 1177 23280 1221 23314
rect 1255 23280 1297 23314
rect 1177 23242 1297 23280
rect 1177 23208 1221 23242
rect 1255 23208 1297 23242
rect 1177 23170 1297 23208
rect 1177 23136 1221 23170
rect 1255 23136 1297 23170
rect 1177 23098 1297 23136
rect 1177 23064 1221 23098
rect 1255 23064 1297 23098
rect 1177 23026 1297 23064
rect 1177 22992 1221 23026
rect 1255 22992 1297 23026
rect 1177 22954 1297 22992
rect 1177 22920 1221 22954
rect 1255 22920 1297 22954
rect 1177 22882 1297 22920
rect 1177 22848 1221 22882
rect 1255 22848 1297 22882
rect 1177 22810 1297 22848
rect 1177 22776 1221 22810
rect 1255 22776 1297 22810
rect 1177 22738 1297 22776
rect 1177 22704 1221 22738
rect 1255 22704 1297 22738
rect 1177 22666 1297 22704
rect 1177 22632 1221 22666
rect 1255 22632 1297 22666
rect 1177 22594 1297 22632
rect 1177 22560 1221 22594
rect 1255 22560 1297 22594
rect 1177 22522 1297 22560
rect 1177 22488 1221 22522
rect 1255 22488 1297 22522
rect 1177 22450 1297 22488
rect 1177 22416 1221 22450
rect 1255 22416 1297 22450
rect 1177 22378 1297 22416
rect 1177 22344 1221 22378
rect 1255 22344 1297 22378
rect 1177 22306 1297 22344
rect 1177 22272 1221 22306
rect 1255 22272 1297 22306
rect 1177 22234 1297 22272
rect 1177 22200 1221 22234
rect 1255 22200 1297 22234
rect 1177 22162 1297 22200
rect 1177 22128 1221 22162
rect 1255 22128 1297 22162
rect 1177 22090 1297 22128
rect 1177 22056 1221 22090
rect 1255 22056 1297 22090
rect 1177 22018 1297 22056
rect 1177 21984 1221 22018
rect 1255 21984 1297 22018
rect 1177 21946 1297 21984
rect 1177 21912 1221 21946
rect 1255 21912 1297 21946
rect 1177 21874 1297 21912
rect 1177 21840 1221 21874
rect 1255 21840 1297 21874
rect 1177 21802 1297 21840
rect 1177 21768 1221 21802
rect 1255 21768 1297 21802
rect 1177 21730 1297 21768
rect 1177 21696 1221 21730
rect 1255 21696 1297 21730
rect 1177 21658 1297 21696
rect 1177 21624 1221 21658
rect 1255 21624 1297 21658
rect 1177 21586 1297 21624
rect 1177 21552 1221 21586
rect 1255 21552 1297 21586
rect 1177 21514 1297 21552
rect 1177 21480 1221 21514
rect 1255 21480 1297 21514
rect 1177 21442 1297 21480
rect 1177 21408 1221 21442
rect 1255 21408 1297 21442
rect 1177 21370 1297 21408
rect 1177 21336 1221 21370
rect 1255 21336 1297 21370
rect 1177 21298 1297 21336
rect 1177 21264 1221 21298
rect 1255 21264 1297 21298
rect 1177 21226 1297 21264
rect 1177 21192 1221 21226
rect 1255 21192 1297 21226
rect 1177 21154 1297 21192
rect 1177 21120 1221 21154
rect 1255 21120 1297 21154
rect 1177 21082 1297 21120
rect 1177 21048 1221 21082
rect 1255 21048 1297 21082
rect 1177 21010 1297 21048
rect 1177 20976 1221 21010
rect 1255 20976 1297 21010
rect 1177 20938 1297 20976
rect 1177 20904 1221 20938
rect 1255 20904 1297 20938
rect 1177 20866 1297 20904
rect 1177 20832 1221 20866
rect 1255 20832 1297 20866
rect 1177 20794 1297 20832
rect 1177 20760 1221 20794
rect 1255 20760 1297 20794
rect 1177 20722 1297 20760
rect 1177 20688 1221 20722
rect 1255 20688 1297 20722
rect 1177 20650 1297 20688
rect 1177 20616 1221 20650
rect 1255 20616 1297 20650
rect 1177 20578 1297 20616
rect 1177 20544 1221 20578
rect 1255 20544 1297 20578
rect 1177 20506 1297 20544
rect 1177 20472 1221 20506
rect 1255 20472 1297 20506
rect 1177 20434 1297 20472
rect 1177 20400 1221 20434
rect 1255 20400 1297 20434
rect 1177 20362 1297 20400
rect 1177 20328 1221 20362
rect 1255 20328 1297 20362
rect 1177 20290 1297 20328
rect 1177 20256 1221 20290
rect 1255 20256 1297 20290
rect 1177 20218 1297 20256
rect 1177 20184 1221 20218
rect 1255 20184 1297 20218
rect 1177 20146 1297 20184
rect 1177 20112 1221 20146
rect 1255 20112 1297 20146
rect 1177 20074 1297 20112
rect 1177 20040 1221 20074
rect 1255 20040 1297 20074
rect 1177 20002 1297 20040
rect 1177 19968 1221 20002
rect 1255 19968 1297 20002
rect 1177 19930 1297 19968
rect 1177 19896 1221 19930
rect 1255 19896 1297 19930
rect 1177 19858 1297 19896
rect 1177 19824 1221 19858
rect 1255 19824 1297 19858
rect 1177 19786 1297 19824
rect 1177 19752 1221 19786
rect 1255 19752 1297 19786
rect 1177 19714 1297 19752
rect 1177 19680 1221 19714
rect 1255 19680 1297 19714
rect 1177 19642 1297 19680
rect 1177 19608 1221 19642
rect 1255 19608 1297 19642
rect 1177 19570 1297 19608
rect 1177 19536 1221 19570
rect 1255 19536 1297 19570
rect 1177 19498 1297 19536
rect 1177 19464 1221 19498
rect 1255 19464 1297 19498
rect 1177 19426 1297 19464
rect 1177 19392 1221 19426
rect 1255 19392 1297 19426
rect 1177 19354 1297 19392
rect 1177 19320 1221 19354
rect 1255 19320 1297 19354
rect 1177 19282 1297 19320
rect 1177 19248 1221 19282
rect 1255 19248 1297 19282
rect 1177 19210 1297 19248
rect 1177 19176 1221 19210
rect 1255 19176 1297 19210
rect 1177 19138 1297 19176
rect 1177 19104 1221 19138
rect 1255 19104 1297 19138
rect 1177 19066 1297 19104
rect 1177 19032 1221 19066
rect 1255 19032 1297 19066
rect 1177 18994 1297 19032
rect 1177 18960 1221 18994
rect 1255 18960 1297 18994
rect 1177 18922 1297 18960
rect 1177 18888 1221 18922
rect 1255 18888 1297 18922
rect 1177 18850 1297 18888
rect 1177 18816 1221 18850
rect 1255 18816 1297 18850
rect 1177 18778 1297 18816
rect 1177 18744 1221 18778
rect 1255 18744 1297 18778
rect 1177 18706 1297 18744
rect 1177 18672 1221 18706
rect 1255 18672 1297 18706
rect 1177 18634 1297 18672
rect 1177 18600 1221 18634
rect 1255 18600 1297 18634
rect 1177 18562 1297 18600
rect 1177 18528 1221 18562
rect 1255 18528 1297 18562
rect 1177 18490 1297 18528
rect 1177 18456 1221 18490
rect 1255 18456 1297 18490
rect 1177 18418 1297 18456
rect 1177 18384 1221 18418
rect 1255 18384 1297 18418
rect 1177 18346 1297 18384
rect 1177 18312 1221 18346
rect 1255 18312 1297 18346
rect 1177 18274 1297 18312
rect 1177 18240 1221 18274
rect 1255 18240 1297 18274
rect 1177 18202 1297 18240
rect 1177 18168 1221 18202
rect 1255 18168 1297 18202
rect 1177 18130 1297 18168
rect 1177 18096 1221 18130
rect 1255 18096 1297 18130
rect 1177 18058 1297 18096
rect 1177 18024 1221 18058
rect 1255 18024 1297 18058
rect 1177 17986 1297 18024
rect 1177 17952 1221 17986
rect 1255 17952 1297 17986
rect 1177 17914 1297 17952
rect 1177 17880 1221 17914
rect 1255 17880 1297 17914
rect 1177 17842 1297 17880
rect 1177 17808 1221 17842
rect 1255 17808 1297 17842
rect 1177 17770 1297 17808
rect 1177 17736 1221 17770
rect 1255 17736 1297 17770
rect 1177 17698 1297 17736
rect 1177 17664 1221 17698
rect 1255 17664 1297 17698
rect 1177 17626 1297 17664
rect 1177 17592 1221 17626
rect 1255 17592 1297 17626
rect 1177 17554 1297 17592
rect 1177 17520 1221 17554
rect 1255 17520 1297 17554
rect 1177 17482 1297 17520
rect 1177 17448 1221 17482
rect 1255 17448 1297 17482
rect 1177 17410 1297 17448
rect 1177 17376 1221 17410
rect 1255 17376 1297 17410
rect 1177 17338 1297 17376
rect 1177 17304 1221 17338
rect 1255 17304 1297 17338
rect 1177 17266 1297 17304
rect 1177 17232 1221 17266
rect 1255 17232 1297 17266
rect 1177 17194 1297 17232
rect 1177 17160 1221 17194
rect 1255 17160 1297 17194
rect 1177 17122 1297 17160
rect 1177 17088 1221 17122
rect 1255 17088 1297 17122
rect 1177 17050 1297 17088
rect 1177 17016 1221 17050
rect 1255 17016 1297 17050
rect 1177 16978 1297 17016
rect 1177 16944 1221 16978
rect 1255 16944 1297 16978
rect 1177 16906 1297 16944
rect 1177 16872 1221 16906
rect 1255 16872 1297 16906
rect 1177 16834 1297 16872
rect 1177 16800 1221 16834
rect 1255 16800 1297 16834
rect 1177 16762 1297 16800
rect 1177 16728 1221 16762
rect 1255 16728 1297 16762
rect 1177 16690 1297 16728
rect 1177 16656 1221 16690
rect 1255 16656 1297 16690
rect 1177 16618 1297 16656
rect 1177 16584 1221 16618
rect 1255 16584 1297 16618
rect 1177 16546 1297 16584
rect 1177 16512 1221 16546
rect 1255 16512 1297 16546
rect 1177 16474 1297 16512
rect 1177 16440 1221 16474
rect 1255 16440 1297 16474
rect 1177 16402 1297 16440
rect 1177 16368 1221 16402
rect 1255 16368 1297 16402
rect 1177 16330 1297 16368
rect 1177 16296 1221 16330
rect 1255 16296 1297 16330
rect 1177 16258 1297 16296
rect 1177 16224 1221 16258
rect 1255 16224 1297 16258
rect 1177 16186 1297 16224
rect 1177 16152 1221 16186
rect 1255 16152 1297 16186
rect 1177 16114 1297 16152
rect 1177 16080 1221 16114
rect 1255 16080 1297 16114
rect 1177 16042 1297 16080
rect 1177 16008 1221 16042
rect 1255 16008 1297 16042
rect 1177 15970 1297 16008
rect 1177 15936 1221 15970
rect 1255 15936 1297 15970
rect 1177 15898 1297 15936
rect 1177 15864 1221 15898
rect 1255 15864 1297 15898
rect 1177 15826 1297 15864
rect 1177 15792 1221 15826
rect 1255 15792 1297 15826
rect 1177 15754 1297 15792
rect 1177 15720 1221 15754
rect 1255 15720 1297 15754
rect 1177 15682 1297 15720
rect 1177 15648 1221 15682
rect 1255 15648 1297 15682
rect 1177 15610 1297 15648
rect 1177 15576 1221 15610
rect 1255 15576 1297 15610
rect 1177 15538 1297 15576
rect 1177 15504 1221 15538
rect 1255 15504 1297 15538
rect 1177 15466 1297 15504
rect 1177 15432 1221 15466
rect 1255 15432 1297 15466
rect 1177 15394 1297 15432
rect 1177 15360 1221 15394
rect 1255 15360 1297 15394
rect 1177 15322 1297 15360
rect 1177 15288 1221 15322
rect 1255 15288 1297 15322
rect 1177 15250 1297 15288
rect 1177 15216 1221 15250
rect 1255 15216 1297 15250
rect 1177 15178 1297 15216
rect 1177 15144 1221 15178
rect 1255 15144 1297 15178
rect 1177 15106 1297 15144
rect 1177 15072 1221 15106
rect 1255 15072 1297 15106
rect 1177 15034 1297 15072
rect 1177 15000 1221 15034
rect 1255 15000 1297 15034
rect 1177 14962 1297 15000
rect 1177 14928 1221 14962
rect 1255 14928 1297 14962
rect 1177 14890 1297 14928
rect 1177 14856 1221 14890
rect 1255 14856 1297 14890
rect 1177 14818 1297 14856
rect 1177 14784 1221 14818
rect 1255 14784 1297 14818
rect 1177 14746 1297 14784
rect 1177 14712 1221 14746
rect 1255 14712 1297 14746
rect 1177 14674 1297 14712
rect 1177 14640 1221 14674
rect 1255 14640 1297 14674
rect 1177 14602 1297 14640
rect 1177 14568 1221 14602
rect 1255 14568 1297 14602
rect 1177 14530 1297 14568
rect 1177 14496 1221 14530
rect 1255 14496 1297 14530
rect 1177 14458 1297 14496
rect 1177 14424 1221 14458
rect 1255 14424 1297 14458
rect 1177 14386 1297 14424
rect 1177 14352 1221 14386
rect 1255 14352 1297 14386
rect 1177 14314 1297 14352
rect 1177 14280 1221 14314
rect 1255 14280 1297 14314
rect 1177 14242 1297 14280
rect 1177 14208 1221 14242
rect 1255 14208 1297 14242
rect 1177 14170 1297 14208
rect 1177 14136 1221 14170
rect 1255 14136 1297 14170
rect 1177 14098 1297 14136
rect 1177 14064 1221 14098
rect 1255 14064 1297 14098
rect 1177 14026 1297 14064
rect 1177 13992 1221 14026
rect 1255 13992 1297 14026
rect 1177 13954 1297 13992
rect 1177 13920 1221 13954
rect 1255 13920 1297 13954
rect 1177 13882 1297 13920
rect 1177 13848 1221 13882
rect 1255 13848 1297 13882
rect 1177 13810 1297 13848
rect 1177 13776 1221 13810
rect 1255 13776 1297 13810
rect 1177 13738 1297 13776
rect 1177 13704 1221 13738
rect 1255 13704 1297 13738
rect 1177 13666 1297 13704
rect 1177 13632 1221 13666
rect 1255 13632 1297 13666
rect 1177 13594 1297 13632
rect 1177 13560 1221 13594
rect 1255 13560 1297 13594
rect 1177 13522 1297 13560
rect 1177 13488 1221 13522
rect 1255 13488 1297 13522
rect 1177 13450 1297 13488
rect 1177 13416 1221 13450
rect 1255 13416 1297 13450
rect 1177 13378 1297 13416
rect 1177 13344 1221 13378
rect 1255 13344 1297 13378
rect 1177 13306 1297 13344
rect 1177 13272 1221 13306
rect 1255 13272 1297 13306
rect 1177 13234 1297 13272
rect 1177 13200 1221 13234
rect 1255 13200 1297 13234
rect 1177 13162 1297 13200
rect 1177 13128 1221 13162
rect 1255 13128 1297 13162
rect 1177 13090 1297 13128
rect 1177 13056 1221 13090
rect 1255 13056 1297 13090
rect 1177 13018 1297 13056
rect 1177 12984 1221 13018
rect 1255 12984 1297 13018
rect 1177 12946 1297 12984
rect 1177 12912 1221 12946
rect 1255 12912 1297 12946
rect 1177 12874 1297 12912
rect 1177 12840 1221 12874
rect 1255 12840 1297 12874
rect 1177 12802 1297 12840
rect 1177 12768 1221 12802
rect 1255 12768 1297 12802
rect 1177 12730 1297 12768
rect 1177 12696 1221 12730
rect 1255 12696 1297 12730
rect 1177 12658 1297 12696
rect 1177 12624 1221 12658
rect 1255 12624 1297 12658
rect 1177 12586 1297 12624
rect 1177 12552 1221 12586
rect 1255 12552 1297 12586
rect 1177 12514 1297 12552
rect 1177 12480 1221 12514
rect 1255 12480 1297 12514
rect 1177 12442 1297 12480
rect 1177 12408 1221 12442
rect 1255 12408 1297 12442
rect 1177 12370 1297 12408
rect 1177 12336 1221 12370
rect 1255 12336 1297 12370
rect 1177 12298 1297 12336
rect 1177 12264 1221 12298
rect 1255 12264 1297 12298
rect 1177 12226 1297 12264
rect 1177 12192 1221 12226
rect 1255 12192 1297 12226
rect 1177 12154 1297 12192
rect 1177 12120 1221 12154
rect 1255 12120 1297 12154
rect 1177 12082 1297 12120
rect 1177 12048 1221 12082
rect 1255 12048 1297 12082
rect 1177 12010 1297 12048
rect 1177 11976 1221 12010
rect 1255 11976 1297 12010
rect 1177 11938 1297 11976
rect 1177 11904 1221 11938
rect 1255 11904 1297 11938
rect 1177 11866 1297 11904
rect 1177 11832 1221 11866
rect 1255 11832 1297 11866
rect 1177 11794 1297 11832
rect 1177 11760 1221 11794
rect 1255 11760 1297 11794
rect 1177 11722 1297 11760
rect 1177 11688 1221 11722
rect 1255 11688 1297 11722
rect 1177 11650 1297 11688
rect 1177 11616 1221 11650
rect 1255 11616 1297 11650
rect 1177 11578 1297 11616
rect 1177 11544 1221 11578
rect 1255 11544 1297 11578
rect 1177 11506 1297 11544
rect 1177 11472 1221 11506
rect 1255 11472 1297 11506
rect 1177 11434 1297 11472
rect 1177 11400 1221 11434
rect 1255 11400 1297 11434
rect 1177 11362 1297 11400
rect 1177 11328 1221 11362
rect 1255 11328 1297 11362
rect 1177 11290 1297 11328
rect 1177 11256 1221 11290
rect 1255 11256 1297 11290
rect 1177 11218 1297 11256
rect 1177 11184 1221 11218
rect 1255 11184 1297 11218
rect 1177 11146 1297 11184
rect 1177 11112 1221 11146
rect 1255 11112 1297 11146
rect 1177 11074 1297 11112
rect 1177 11040 1221 11074
rect 1255 11040 1297 11074
rect 1177 11002 1297 11040
rect 1177 10968 1221 11002
rect 1255 10968 1297 11002
rect 1177 10930 1297 10968
rect 1177 10896 1221 10930
rect 1255 10896 1297 10930
rect 1177 10858 1297 10896
rect 1177 10824 1221 10858
rect 1255 10824 1297 10858
rect 1177 10786 1297 10824
rect 13697 34478 13817 34564
rect 13697 34444 13739 34478
rect 13773 34444 13817 34478
rect 13697 34406 13817 34444
rect 13697 34372 13739 34406
rect 13773 34372 13817 34406
rect 13697 34334 13817 34372
rect 13697 34300 13739 34334
rect 13773 34300 13817 34334
rect 13697 34262 13817 34300
rect 13697 34228 13739 34262
rect 13773 34228 13817 34262
rect 13697 34190 13817 34228
rect 13697 34156 13739 34190
rect 13773 34156 13817 34190
rect 13697 34118 13817 34156
rect 13697 34084 13739 34118
rect 13773 34084 13817 34118
rect 13697 34046 13817 34084
rect 13697 34012 13739 34046
rect 13773 34012 13817 34046
rect 13697 33974 13817 34012
rect 13697 33940 13739 33974
rect 13773 33940 13817 33974
rect 13697 33902 13817 33940
rect 13697 33868 13739 33902
rect 13773 33868 13817 33902
rect 13697 33830 13817 33868
rect 13697 33796 13739 33830
rect 13773 33796 13817 33830
rect 13697 33758 13817 33796
rect 13697 33724 13739 33758
rect 13773 33724 13817 33758
rect 13697 33686 13817 33724
rect 13697 33652 13739 33686
rect 13773 33652 13817 33686
rect 13697 33614 13817 33652
rect 13697 33580 13739 33614
rect 13773 33580 13817 33614
rect 13697 33542 13817 33580
rect 13697 33508 13739 33542
rect 13773 33508 13817 33542
rect 13697 33470 13817 33508
rect 13697 33436 13739 33470
rect 13773 33436 13817 33470
rect 13697 33398 13817 33436
rect 13697 33364 13739 33398
rect 13773 33364 13817 33398
rect 13697 33326 13817 33364
rect 13697 33292 13739 33326
rect 13773 33292 13817 33326
rect 13697 33254 13817 33292
rect 13697 33220 13739 33254
rect 13773 33220 13817 33254
rect 13697 33182 13817 33220
rect 13697 33148 13739 33182
rect 13773 33148 13817 33182
rect 13697 33110 13817 33148
rect 13697 33076 13739 33110
rect 13773 33076 13817 33110
rect 13697 33038 13817 33076
rect 13697 33004 13739 33038
rect 13773 33004 13817 33038
rect 13697 32966 13817 33004
rect 13697 32932 13739 32966
rect 13773 32932 13817 32966
rect 13697 32894 13817 32932
rect 13697 32860 13739 32894
rect 13773 32860 13817 32894
rect 13697 32822 13817 32860
rect 13697 32788 13739 32822
rect 13773 32788 13817 32822
rect 13697 32750 13817 32788
rect 13697 32716 13739 32750
rect 13773 32716 13817 32750
rect 13697 32678 13817 32716
rect 13697 32644 13739 32678
rect 13773 32644 13817 32678
rect 13697 32606 13817 32644
rect 13697 32572 13739 32606
rect 13773 32572 13817 32606
rect 13697 32534 13817 32572
rect 13697 32500 13739 32534
rect 13773 32500 13817 32534
rect 13697 32462 13817 32500
rect 13697 32428 13739 32462
rect 13773 32428 13817 32462
rect 13697 32390 13817 32428
rect 13697 32356 13739 32390
rect 13773 32356 13817 32390
rect 13697 32318 13817 32356
rect 13697 32284 13739 32318
rect 13773 32284 13817 32318
rect 13697 32246 13817 32284
rect 13697 32212 13739 32246
rect 13773 32212 13817 32246
rect 13697 32174 13817 32212
rect 13697 32140 13739 32174
rect 13773 32140 13817 32174
rect 13697 32102 13817 32140
rect 13697 32068 13739 32102
rect 13773 32068 13817 32102
rect 13697 32030 13817 32068
rect 13697 31996 13739 32030
rect 13773 31996 13817 32030
rect 13697 31958 13817 31996
rect 13697 31924 13739 31958
rect 13773 31924 13817 31958
rect 13697 31886 13817 31924
rect 13697 31852 13739 31886
rect 13773 31852 13817 31886
rect 13697 31814 13817 31852
rect 13697 31780 13739 31814
rect 13773 31780 13817 31814
rect 13697 31742 13817 31780
rect 13697 31708 13739 31742
rect 13773 31708 13817 31742
rect 13697 31670 13817 31708
rect 13697 31636 13739 31670
rect 13773 31636 13817 31670
rect 13697 31598 13817 31636
rect 13697 31564 13739 31598
rect 13773 31564 13817 31598
rect 13697 31526 13817 31564
rect 13697 31492 13739 31526
rect 13773 31492 13817 31526
rect 13697 31454 13817 31492
rect 13697 31420 13739 31454
rect 13773 31420 13817 31454
rect 13697 31382 13817 31420
rect 13697 31348 13739 31382
rect 13773 31348 13817 31382
rect 13697 31310 13817 31348
rect 13697 31276 13739 31310
rect 13773 31276 13817 31310
rect 13697 31238 13817 31276
rect 13697 31204 13739 31238
rect 13773 31204 13817 31238
rect 13697 31166 13817 31204
rect 13697 31132 13739 31166
rect 13773 31132 13817 31166
rect 13697 31094 13817 31132
rect 13697 31060 13739 31094
rect 13773 31060 13817 31094
rect 13697 31022 13817 31060
rect 13697 30988 13739 31022
rect 13773 30988 13817 31022
rect 13697 30950 13817 30988
rect 13697 30916 13739 30950
rect 13773 30916 13817 30950
rect 13697 30878 13817 30916
rect 13697 30844 13739 30878
rect 13773 30844 13817 30878
rect 13697 30806 13817 30844
rect 13697 30772 13739 30806
rect 13773 30772 13817 30806
rect 13697 30734 13817 30772
rect 13697 30700 13739 30734
rect 13773 30700 13817 30734
rect 13697 30662 13817 30700
rect 13697 30628 13739 30662
rect 13773 30628 13817 30662
rect 13697 30590 13817 30628
rect 13697 30556 13739 30590
rect 13773 30556 13817 30590
rect 13697 30518 13817 30556
rect 13697 30484 13739 30518
rect 13773 30484 13817 30518
rect 13697 30446 13817 30484
rect 13697 30412 13739 30446
rect 13773 30412 13817 30446
rect 13697 30374 13817 30412
rect 13697 30340 13739 30374
rect 13773 30340 13817 30374
rect 13697 30302 13817 30340
rect 13697 30268 13739 30302
rect 13773 30268 13817 30302
rect 13697 30230 13817 30268
rect 13697 30196 13739 30230
rect 13773 30196 13817 30230
rect 13697 30158 13817 30196
rect 13697 30124 13739 30158
rect 13773 30124 13817 30158
rect 13697 30086 13817 30124
rect 13697 30052 13739 30086
rect 13773 30052 13817 30086
rect 13697 30014 13817 30052
rect 13697 29980 13739 30014
rect 13773 29980 13817 30014
rect 13697 29942 13817 29980
rect 13697 29908 13739 29942
rect 13773 29908 13817 29942
rect 13697 29870 13817 29908
rect 13697 29836 13739 29870
rect 13773 29836 13817 29870
rect 13697 29798 13817 29836
rect 13697 29764 13739 29798
rect 13773 29764 13817 29798
rect 13697 29726 13817 29764
rect 13697 29692 13739 29726
rect 13773 29692 13817 29726
rect 13697 29654 13817 29692
rect 13697 29620 13739 29654
rect 13773 29620 13817 29654
rect 13697 29582 13817 29620
rect 13697 29548 13739 29582
rect 13773 29548 13817 29582
rect 13697 29510 13817 29548
rect 13697 29476 13739 29510
rect 13773 29476 13817 29510
rect 13697 29438 13817 29476
rect 13697 29404 13739 29438
rect 13773 29404 13817 29438
rect 13697 29366 13817 29404
rect 13697 29332 13739 29366
rect 13773 29332 13817 29366
rect 13697 29294 13817 29332
rect 13697 29260 13739 29294
rect 13773 29260 13817 29294
rect 13697 29222 13817 29260
rect 13697 29188 13739 29222
rect 13773 29188 13817 29222
rect 13697 29150 13817 29188
rect 13697 29116 13739 29150
rect 13773 29116 13817 29150
rect 13697 29078 13817 29116
rect 13697 29044 13739 29078
rect 13773 29044 13817 29078
rect 13697 29006 13817 29044
rect 13697 28972 13739 29006
rect 13773 28972 13817 29006
rect 13697 28934 13817 28972
rect 13697 28900 13739 28934
rect 13773 28900 13817 28934
rect 13697 28862 13817 28900
rect 13697 28828 13739 28862
rect 13773 28828 13817 28862
rect 13697 28790 13817 28828
rect 13697 28756 13739 28790
rect 13773 28756 13817 28790
rect 13697 28718 13817 28756
rect 13697 28684 13739 28718
rect 13773 28684 13817 28718
rect 13697 28646 13817 28684
rect 13697 28612 13739 28646
rect 13773 28612 13817 28646
rect 13697 28574 13817 28612
rect 13697 28540 13739 28574
rect 13773 28540 13817 28574
rect 13697 28502 13817 28540
rect 13697 28468 13739 28502
rect 13773 28468 13817 28502
rect 13697 28430 13817 28468
rect 13697 28396 13739 28430
rect 13773 28396 13817 28430
rect 13697 28358 13817 28396
rect 13697 28324 13739 28358
rect 13773 28324 13817 28358
rect 13697 28286 13817 28324
rect 13697 28252 13739 28286
rect 13773 28252 13817 28286
rect 13697 28214 13817 28252
rect 13697 28180 13739 28214
rect 13773 28180 13817 28214
rect 13697 28142 13817 28180
rect 13697 28108 13739 28142
rect 13773 28108 13817 28142
rect 13697 28070 13817 28108
rect 13697 28036 13739 28070
rect 13773 28036 13817 28070
rect 13697 27998 13817 28036
rect 13697 27964 13739 27998
rect 13773 27964 13817 27998
rect 13697 27926 13817 27964
rect 13697 27892 13739 27926
rect 13773 27892 13817 27926
rect 13697 27854 13817 27892
rect 13697 27820 13739 27854
rect 13773 27820 13817 27854
rect 13697 27782 13817 27820
rect 13697 27748 13739 27782
rect 13773 27748 13817 27782
rect 13697 27710 13817 27748
rect 13697 27676 13739 27710
rect 13773 27676 13817 27710
rect 13697 27638 13817 27676
rect 13697 27604 13739 27638
rect 13773 27604 13817 27638
rect 13697 27566 13817 27604
rect 13697 27532 13739 27566
rect 13773 27532 13817 27566
rect 13697 27494 13817 27532
rect 13697 27460 13739 27494
rect 13773 27460 13817 27494
rect 13697 27422 13817 27460
rect 13697 27388 13739 27422
rect 13773 27388 13817 27422
rect 13697 27350 13817 27388
rect 13697 27316 13739 27350
rect 13773 27316 13817 27350
rect 13697 27278 13817 27316
rect 13697 27244 13739 27278
rect 13773 27244 13817 27278
rect 13697 27206 13817 27244
rect 13697 27172 13739 27206
rect 13773 27172 13817 27206
rect 13697 27134 13817 27172
rect 13697 27100 13739 27134
rect 13773 27100 13817 27134
rect 13697 27062 13817 27100
rect 13697 27028 13739 27062
rect 13773 27028 13817 27062
rect 13697 26990 13817 27028
rect 13697 26956 13739 26990
rect 13773 26956 13817 26990
rect 13697 26918 13817 26956
rect 13697 26884 13739 26918
rect 13773 26884 13817 26918
rect 13697 26846 13817 26884
rect 13697 26812 13739 26846
rect 13773 26812 13817 26846
rect 13697 26774 13817 26812
rect 13697 26740 13739 26774
rect 13773 26740 13817 26774
rect 13697 26702 13817 26740
rect 13697 26668 13739 26702
rect 13773 26668 13817 26702
rect 13697 26630 13817 26668
rect 13697 26596 13739 26630
rect 13773 26596 13817 26630
rect 13697 26558 13817 26596
rect 13697 26524 13739 26558
rect 13773 26524 13817 26558
rect 13697 26486 13817 26524
rect 13697 26452 13739 26486
rect 13773 26452 13817 26486
rect 13697 26414 13817 26452
rect 13697 26380 13739 26414
rect 13773 26380 13817 26414
rect 13697 26342 13817 26380
rect 13697 26308 13739 26342
rect 13773 26308 13817 26342
rect 13697 26270 13817 26308
rect 13697 26236 13739 26270
rect 13773 26236 13817 26270
rect 13697 26198 13817 26236
rect 13697 26164 13739 26198
rect 13773 26164 13817 26198
rect 13697 26126 13817 26164
rect 13697 26092 13739 26126
rect 13773 26092 13817 26126
rect 13697 26054 13817 26092
rect 13697 26020 13739 26054
rect 13773 26020 13817 26054
rect 13697 25982 13817 26020
rect 13697 25948 13739 25982
rect 13773 25948 13817 25982
rect 13697 25910 13817 25948
rect 13697 25876 13739 25910
rect 13773 25876 13817 25910
rect 13697 25838 13817 25876
rect 13697 25804 13739 25838
rect 13773 25804 13817 25838
rect 13697 25766 13817 25804
rect 13697 25732 13739 25766
rect 13773 25732 13817 25766
rect 13697 25694 13817 25732
rect 13697 25660 13739 25694
rect 13773 25660 13817 25694
rect 13697 25622 13817 25660
rect 13697 25588 13739 25622
rect 13773 25588 13817 25622
rect 13697 25550 13817 25588
rect 13697 25516 13739 25550
rect 13773 25516 13817 25550
rect 13697 25478 13817 25516
rect 13697 25444 13739 25478
rect 13773 25444 13817 25478
rect 13697 25406 13817 25444
rect 13697 25372 13739 25406
rect 13773 25372 13817 25406
rect 13697 25334 13817 25372
rect 13697 25300 13739 25334
rect 13773 25300 13817 25334
rect 13697 25262 13817 25300
rect 13697 25228 13739 25262
rect 13773 25228 13817 25262
rect 13697 25190 13817 25228
rect 13697 25156 13739 25190
rect 13773 25156 13817 25190
rect 13697 25118 13817 25156
rect 13697 25084 13739 25118
rect 13773 25084 13817 25118
rect 13697 25046 13817 25084
rect 13697 25012 13739 25046
rect 13773 25012 13817 25046
rect 13697 24974 13817 25012
rect 13697 24940 13739 24974
rect 13773 24940 13817 24974
rect 13697 24902 13817 24940
rect 13697 24868 13739 24902
rect 13773 24868 13817 24902
rect 13697 24830 13817 24868
rect 13697 24796 13739 24830
rect 13773 24796 13817 24830
rect 13697 24758 13817 24796
rect 13697 24724 13739 24758
rect 13773 24724 13817 24758
rect 13697 24686 13817 24724
rect 13697 24652 13739 24686
rect 13773 24652 13817 24686
rect 13697 24614 13817 24652
rect 13697 24580 13739 24614
rect 13773 24580 13817 24614
rect 13697 24542 13817 24580
rect 13697 24508 13739 24542
rect 13773 24508 13817 24542
rect 13697 24470 13817 24508
rect 13697 24436 13739 24470
rect 13773 24436 13817 24470
rect 13697 24398 13817 24436
rect 13697 24364 13739 24398
rect 13773 24364 13817 24398
rect 13697 24326 13817 24364
rect 13697 24292 13739 24326
rect 13773 24292 13817 24326
rect 13697 24254 13817 24292
rect 13697 24220 13739 24254
rect 13773 24220 13817 24254
rect 13697 24182 13817 24220
rect 13697 24148 13739 24182
rect 13773 24148 13817 24182
rect 13697 24110 13817 24148
rect 13697 24076 13739 24110
rect 13773 24076 13817 24110
rect 13697 24038 13817 24076
rect 13697 24004 13739 24038
rect 13773 24004 13817 24038
rect 13697 23966 13817 24004
rect 13697 23932 13739 23966
rect 13773 23932 13817 23966
rect 13697 23894 13817 23932
rect 13697 23860 13739 23894
rect 13773 23860 13817 23894
rect 13697 23822 13817 23860
rect 13697 23788 13739 23822
rect 13773 23788 13817 23822
rect 13697 23750 13817 23788
rect 13697 23716 13739 23750
rect 13773 23716 13817 23750
rect 13697 23678 13817 23716
rect 13697 23644 13739 23678
rect 13773 23644 13817 23678
rect 13697 23606 13817 23644
rect 13697 23572 13739 23606
rect 13773 23572 13817 23606
rect 13697 23534 13817 23572
rect 13697 23500 13739 23534
rect 13773 23500 13817 23534
rect 13697 23462 13817 23500
rect 13697 23428 13739 23462
rect 13773 23428 13817 23462
rect 13697 23390 13817 23428
rect 13697 23356 13739 23390
rect 13773 23356 13817 23390
rect 13697 23318 13817 23356
rect 13697 23284 13739 23318
rect 13773 23284 13817 23318
rect 13697 23246 13817 23284
rect 13697 23212 13739 23246
rect 13773 23212 13817 23246
rect 13697 23174 13817 23212
rect 13697 23140 13739 23174
rect 13773 23140 13817 23174
rect 13697 23102 13817 23140
rect 13697 23068 13739 23102
rect 13773 23068 13817 23102
rect 13697 23030 13817 23068
rect 13697 22996 13739 23030
rect 13773 22996 13817 23030
rect 13697 22958 13817 22996
rect 13697 22924 13739 22958
rect 13773 22924 13817 22958
rect 13697 22886 13817 22924
rect 13697 22852 13739 22886
rect 13773 22852 13817 22886
rect 13697 22814 13817 22852
rect 13697 22780 13739 22814
rect 13773 22780 13817 22814
rect 13697 22742 13817 22780
rect 13697 22708 13739 22742
rect 13773 22708 13817 22742
rect 13697 22670 13817 22708
rect 13697 22636 13739 22670
rect 13773 22636 13817 22670
rect 13697 22598 13817 22636
rect 13697 22564 13739 22598
rect 13773 22564 13817 22598
rect 13697 22526 13817 22564
rect 13697 22492 13739 22526
rect 13773 22492 13817 22526
rect 13697 22454 13817 22492
rect 13697 22420 13739 22454
rect 13773 22420 13817 22454
rect 13697 22382 13817 22420
rect 13697 22348 13739 22382
rect 13773 22348 13817 22382
rect 13697 22310 13817 22348
rect 13697 22276 13739 22310
rect 13773 22276 13817 22310
rect 13697 22238 13817 22276
rect 13697 22204 13739 22238
rect 13773 22204 13817 22238
rect 13697 22166 13817 22204
rect 13697 22132 13739 22166
rect 13773 22132 13817 22166
rect 13697 22094 13817 22132
rect 13697 22060 13739 22094
rect 13773 22060 13817 22094
rect 13697 22022 13817 22060
rect 13697 21988 13739 22022
rect 13773 21988 13817 22022
rect 13697 21950 13817 21988
rect 13697 21916 13739 21950
rect 13773 21916 13817 21950
rect 13697 21878 13817 21916
rect 13697 21844 13739 21878
rect 13773 21844 13817 21878
rect 13697 21806 13817 21844
rect 13697 21772 13739 21806
rect 13773 21772 13817 21806
rect 13697 21734 13817 21772
rect 13697 21700 13739 21734
rect 13773 21700 13817 21734
rect 13697 21662 13817 21700
rect 13697 21628 13739 21662
rect 13773 21628 13817 21662
rect 13697 21590 13817 21628
rect 13697 21556 13739 21590
rect 13773 21556 13817 21590
rect 13697 21518 13817 21556
rect 13697 21484 13739 21518
rect 13773 21484 13817 21518
rect 13697 21446 13817 21484
rect 13697 21412 13739 21446
rect 13773 21412 13817 21446
rect 13697 21374 13817 21412
rect 13697 21340 13739 21374
rect 13773 21340 13817 21374
rect 13697 21302 13817 21340
rect 13697 21268 13739 21302
rect 13773 21268 13817 21302
rect 13697 21230 13817 21268
rect 13697 21196 13739 21230
rect 13773 21196 13817 21230
rect 13697 21158 13817 21196
rect 13697 21124 13739 21158
rect 13773 21124 13817 21158
rect 13697 21086 13817 21124
rect 13697 21052 13739 21086
rect 13773 21052 13817 21086
rect 13697 21014 13817 21052
rect 13697 20980 13739 21014
rect 13773 20980 13817 21014
rect 13697 20942 13817 20980
rect 13697 20908 13739 20942
rect 13773 20908 13817 20942
rect 13697 20870 13817 20908
rect 13697 20836 13739 20870
rect 13773 20836 13817 20870
rect 13697 20798 13817 20836
rect 13697 20764 13739 20798
rect 13773 20764 13817 20798
rect 13697 20726 13817 20764
rect 13697 20692 13739 20726
rect 13773 20692 13817 20726
rect 13697 20654 13817 20692
rect 13697 20620 13739 20654
rect 13773 20620 13817 20654
rect 13697 20582 13817 20620
rect 13697 20548 13739 20582
rect 13773 20548 13817 20582
rect 13697 20510 13817 20548
rect 13697 20476 13739 20510
rect 13773 20476 13817 20510
rect 13697 20438 13817 20476
rect 13697 20404 13739 20438
rect 13773 20404 13817 20438
rect 13697 20366 13817 20404
rect 13697 20332 13739 20366
rect 13773 20332 13817 20366
rect 13697 20294 13817 20332
rect 13697 20260 13739 20294
rect 13773 20260 13817 20294
rect 13697 20222 13817 20260
rect 13697 20188 13739 20222
rect 13773 20188 13817 20222
rect 13697 20150 13817 20188
rect 13697 20116 13739 20150
rect 13773 20116 13817 20150
rect 13697 20078 13817 20116
rect 13697 20044 13739 20078
rect 13773 20044 13817 20078
rect 13697 20006 13817 20044
rect 13697 19972 13739 20006
rect 13773 19972 13817 20006
rect 13697 19934 13817 19972
rect 13697 19900 13739 19934
rect 13773 19900 13817 19934
rect 13697 19862 13817 19900
rect 13697 19828 13739 19862
rect 13773 19828 13817 19862
rect 13697 19790 13817 19828
rect 13697 19756 13739 19790
rect 13773 19756 13817 19790
rect 13697 19718 13817 19756
rect 13697 19684 13739 19718
rect 13773 19684 13817 19718
rect 13697 19646 13817 19684
rect 13697 19612 13739 19646
rect 13773 19612 13817 19646
rect 13697 19574 13817 19612
rect 13697 19540 13739 19574
rect 13773 19540 13817 19574
rect 13697 19502 13817 19540
rect 13697 19468 13739 19502
rect 13773 19468 13817 19502
rect 13697 19430 13817 19468
rect 13697 19396 13739 19430
rect 13773 19396 13817 19430
rect 13697 19358 13817 19396
rect 13697 19324 13739 19358
rect 13773 19324 13817 19358
rect 13697 19286 13817 19324
rect 13697 19252 13739 19286
rect 13773 19252 13817 19286
rect 13697 19214 13817 19252
rect 13697 19180 13739 19214
rect 13773 19180 13817 19214
rect 13697 19142 13817 19180
rect 13697 19108 13739 19142
rect 13773 19108 13817 19142
rect 13697 19070 13817 19108
rect 13697 19036 13739 19070
rect 13773 19036 13817 19070
rect 13697 18998 13817 19036
rect 13697 18964 13739 18998
rect 13773 18964 13817 18998
rect 13697 18926 13817 18964
rect 13697 18892 13739 18926
rect 13773 18892 13817 18926
rect 13697 18854 13817 18892
rect 13697 18820 13739 18854
rect 13773 18820 13817 18854
rect 13697 18782 13817 18820
rect 13697 18748 13739 18782
rect 13773 18748 13817 18782
rect 13697 18710 13817 18748
rect 13697 18676 13739 18710
rect 13773 18676 13817 18710
rect 13697 18638 13817 18676
rect 13697 18604 13739 18638
rect 13773 18604 13817 18638
rect 13697 18566 13817 18604
rect 13697 18532 13739 18566
rect 13773 18532 13817 18566
rect 13697 18494 13817 18532
rect 13697 18460 13739 18494
rect 13773 18460 13817 18494
rect 13697 18422 13817 18460
rect 13697 18388 13739 18422
rect 13773 18388 13817 18422
rect 13697 18350 13817 18388
rect 13697 18316 13739 18350
rect 13773 18316 13817 18350
rect 13697 18278 13817 18316
rect 13697 18244 13739 18278
rect 13773 18244 13817 18278
rect 13697 18206 13817 18244
rect 13697 18172 13739 18206
rect 13773 18172 13817 18206
rect 13697 18134 13817 18172
rect 13697 18100 13739 18134
rect 13773 18100 13817 18134
rect 13697 18062 13817 18100
rect 13697 18028 13739 18062
rect 13773 18028 13817 18062
rect 13697 17990 13817 18028
rect 13697 17956 13739 17990
rect 13773 17956 13817 17990
rect 13697 17918 13817 17956
rect 13697 17884 13739 17918
rect 13773 17884 13817 17918
rect 13697 17846 13817 17884
rect 13697 17812 13739 17846
rect 13773 17812 13817 17846
rect 13697 17774 13817 17812
rect 13697 17740 13739 17774
rect 13773 17740 13817 17774
rect 13697 17702 13817 17740
rect 13697 17668 13739 17702
rect 13773 17668 13817 17702
rect 13697 17630 13817 17668
rect 13697 17596 13739 17630
rect 13773 17596 13817 17630
rect 13697 17558 13817 17596
rect 13697 17524 13739 17558
rect 13773 17524 13817 17558
rect 13697 17486 13817 17524
rect 13697 17452 13739 17486
rect 13773 17452 13817 17486
rect 13697 17414 13817 17452
rect 13697 17380 13739 17414
rect 13773 17380 13817 17414
rect 13697 17342 13817 17380
rect 13697 17308 13739 17342
rect 13773 17308 13817 17342
rect 13697 17270 13817 17308
rect 13697 17236 13739 17270
rect 13773 17236 13817 17270
rect 13697 17198 13817 17236
rect 13697 17164 13739 17198
rect 13773 17164 13817 17198
rect 13697 17126 13817 17164
rect 13697 17092 13739 17126
rect 13773 17092 13817 17126
rect 13697 17054 13817 17092
rect 13697 17020 13739 17054
rect 13773 17020 13817 17054
rect 13697 16982 13817 17020
rect 13697 16948 13739 16982
rect 13773 16948 13817 16982
rect 13697 16910 13817 16948
rect 13697 16876 13739 16910
rect 13773 16876 13817 16910
rect 13697 16838 13817 16876
rect 13697 16804 13739 16838
rect 13773 16804 13817 16838
rect 13697 16766 13817 16804
rect 13697 16732 13739 16766
rect 13773 16732 13817 16766
rect 13697 16694 13817 16732
rect 13697 16660 13739 16694
rect 13773 16660 13817 16694
rect 13697 16622 13817 16660
rect 13697 16588 13739 16622
rect 13773 16588 13817 16622
rect 13697 16550 13817 16588
rect 13697 16516 13739 16550
rect 13773 16516 13817 16550
rect 13697 16478 13817 16516
rect 13697 16444 13739 16478
rect 13773 16444 13817 16478
rect 13697 16406 13817 16444
rect 13697 16372 13739 16406
rect 13773 16372 13817 16406
rect 13697 16334 13817 16372
rect 13697 16300 13739 16334
rect 13773 16300 13817 16334
rect 13697 16262 13817 16300
rect 13697 16228 13739 16262
rect 13773 16228 13817 16262
rect 13697 16190 13817 16228
rect 13697 16156 13739 16190
rect 13773 16156 13817 16190
rect 13697 16118 13817 16156
rect 13697 16084 13739 16118
rect 13773 16084 13817 16118
rect 13697 16046 13817 16084
rect 13697 16012 13739 16046
rect 13773 16012 13817 16046
rect 13697 15974 13817 16012
rect 13697 15940 13739 15974
rect 13773 15940 13817 15974
rect 13697 15902 13817 15940
rect 13697 15868 13739 15902
rect 13773 15868 13817 15902
rect 13697 15830 13817 15868
rect 13697 15796 13739 15830
rect 13773 15796 13817 15830
rect 13697 15758 13817 15796
rect 13697 15724 13739 15758
rect 13773 15724 13817 15758
rect 13697 15686 13817 15724
rect 13697 15652 13739 15686
rect 13773 15652 13817 15686
rect 13697 15614 13817 15652
rect 13697 15580 13739 15614
rect 13773 15580 13817 15614
rect 13697 15542 13817 15580
rect 13697 15508 13739 15542
rect 13773 15508 13817 15542
rect 13697 15470 13817 15508
rect 13697 15436 13739 15470
rect 13773 15436 13817 15470
rect 13697 15398 13817 15436
rect 13697 15364 13739 15398
rect 13773 15364 13817 15398
rect 13697 15326 13817 15364
rect 13697 15292 13739 15326
rect 13773 15292 13817 15326
rect 13697 15254 13817 15292
rect 13697 15220 13739 15254
rect 13773 15220 13817 15254
rect 13697 15182 13817 15220
rect 13697 15148 13739 15182
rect 13773 15148 13817 15182
rect 13697 15110 13817 15148
rect 13697 15076 13739 15110
rect 13773 15076 13817 15110
rect 13697 15038 13817 15076
rect 13697 15004 13739 15038
rect 13773 15004 13817 15038
rect 13697 14966 13817 15004
rect 13697 14932 13739 14966
rect 13773 14932 13817 14966
rect 13697 14894 13817 14932
rect 13697 14860 13739 14894
rect 13773 14860 13817 14894
rect 13697 14822 13817 14860
rect 13697 14788 13739 14822
rect 13773 14788 13817 14822
rect 13697 14750 13817 14788
rect 13697 14716 13739 14750
rect 13773 14716 13817 14750
rect 13697 14678 13817 14716
rect 13697 14644 13739 14678
rect 13773 14644 13817 14678
rect 13697 14606 13817 14644
rect 13697 14572 13739 14606
rect 13773 14572 13817 14606
rect 13697 14534 13817 14572
rect 13697 14500 13739 14534
rect 13773 14500 13817 14534
rect 13697 14462 13817 14500
rect 13697 14428 13739 14462
rect 13773 14428 13817 14462
rect 13697 14390 13817 14428
rect 13697 14356 13739 14390
rect 13773 14356 13817 14390
rect 13697 14318 13817 14356
rect 13697 14284 13739 14318
rect 13773 14284 13817 14318
rect 13697 14246 13817 14284
rect 13697 14212 13739 14246
rect 13773 14212 13817 14246
rect 13697 14174 13817 14212
rect 13697 14140 13739 14174
rect 13773 14140 13817 14174
rect 13697 14102 13817 14140
rect 13697 14068 13739 14102
rect 13773 14068 13817 14102
rect 13697 14030 13817 14068
rect 13697 13996 13739 14030
rect 13773 13996 13817 14030
rect 13697 13958 13817 13996
rect 13697 13924 13739 13958
rect 13773 13924 13817 13958
rect 13697 13886 13817 13924
rect 13697 13852 13739 13886
rect 13773 13852 13817 13886
rect 13697 13814 13817 13852
rect 13697 13780 13739 13814
rect 13773 13780 13817 13814
rect 13697 13742 13817 13780
rect 13697 13708 13739 13742
rect 13773 13708 13817 13742
rect 13697 13670 13817 13708
rect 13697 13636 13739 13670
rect 13773 13636 13817 13670
rect 13697 13598 13817 13636
rect 13697 13564 13739 13598
rect 13773 13564 13817 13598
rect 13697 13526 13817 13564
rect 13697 13492 13739 13526
rect 13773 13492 13817 13526
rect 13697 13454 13817 13492
rect 13697 13420 13739 13454
rect 13773 13420 13817 13454
rect 13697 13382 13817 13420
rect 13697 13348 13739 13382
rect 13773 13348 13817 13382
rect 13697 13310 13817 13348
rect 13697 13276 13739 13310
rect 13773 13276 13817 13310
rect 13697 13238 13817 13276
rect 13697 13204 13739 13238
rect 13773 13204 13817 13238
rect 13697 13166 13817 13204
rect 13697 13132 13739 13166
rect 13773 13132 13817 13166
rect 13697 13094 13817 13132
rect 13697 13060 13739 13094
rect 13773 13060 13817 13094
rect 13697 13022 13817 13060
rect 13697 12988 13739 13022
rect 13773 12988 13817 13022
rect 13697 12950 13817 12988
rect 13697 12916 13739 12950
rect 13773 12916 13817 12950
rect 13697 12878 13817 12916
rect 13697 12844 13739 12878
rect 13773 12844 13817 12878
rect 13697 12806 13817 12844
rect 13697 12772 13739 12806
rect 13773 12772 13817 12806
rect 13697 12734 13817 12772
rect 13697 12700 13739 12734
rect 13773 12700 13817 12734
rect 13697 12662 13817 12700
rect 13697 12628 13739 12662
rect 13773 12628 13817 12662
rect 13697 12590 13817 12628
rect 13697 12556 13739 12590
rect 13773 12556 13817 12590
rect 13697 12518 13817 12556
rect 13697 12484 13739 12518
rect 13773 12484 13817 12518
rect 13697 12446 13817 12484
rect 13697 12412 13739 12446
rect 13773 12412 13817 12446
rect 13697 12374 13817 12412
rect 13697 12340 13739 12374
rect 13773 12340 13817 12374
rect 13697 12302 13817 12340
rect 13697 12268 13739 12302
rect 13773 12268 13817 12302
rect 13697 12230 13817 12268
rect 13697 12196 13739 12230
rect 13773 12196 13817 12230
rect 13697 12158 13817 12196
rect 13697 12124 13739 12158
rect 13773 12124 13817 12158
rect 13697 12086 13817 12124
rect 13697 12052 13739 12086
rect 13773 12052 13817 12086
rect 13697 12014 13817 12052
rect 13697 11980 13739 12014
rect 13773 11980 13817 12014
rect 13697 11942 13817 11980
rect 13697 11908 13739 11942
rect 13773 11908 13817 11942
rect 13697 11870 13817 11908
rect 13697 11836 13739 11870
rect 13773 11836 13817 11870
rect 13697 11798 13817 11836
rect 13697 11764 13739 11798
rect 13773 11764 13817 11798
rect 13697 11726 13817 11764
rect 13697 11692 13739 11726
rect 13773 11692 13817 11726
rect 13697 11654 13817 11692
rect 13697 11620 13739 11654
rect 13773 11620 13817 11654
rect 13697 11582 13817 11620
rect 13697 11548 13739 11582
rect 13773 11548 13817 11582
rect 13697 11510 13817 11548
rect 13697 11476 13739 11510
rect 13773 11476 13817 11510
rect 13697 11438 13817 11476
rect 13697 11404 13739 11438
rect 13773 11404 13817 11438
rect 13697 11366 13817 11404
rect 13697 11332 13739 11366
rect 13773 11332 13817 11366
rect 13697 11294 13817 11332
rect 13697 11260 13739 11294
rect 13773 11260 13817 11294
rect 13697 11222 13817 11260
rect 13697 11188 13739 11222
rect 13773 11188 13817 11222
rect 13697 11150 13817 11188
rect 13697 11116 13739 11150
rect 13773 11116 13817 11150
rect 13697 11078 13817 11116
rect 13697 11044 13739 11078
rect 13773 11044 13817 11078
rect 13697 11006 13817 11044
rect 13697 10972 13739 11006
rect 13773 10972 13817 11006
rect 13697 10934 13817 10972
rect 13697 10900 13739 10934
rect 13773 10900 13817 10934
rect 13697 10862 13817 10900
rect 13697 10828 13739 10862
rect 13773 10828 13817 10862
rect 1177 10752 1221 10786
rect 1255 10752 1297 10786
rect 1177 10714 1297 10752
rect 1177 10680 1221 10714
rect 1255 10680 1297 10714
rect 1177 10642 1297 10680
rect 1177 10608 1221 10642
rect 1255 10608 1297 10642
rect 1177 10570 1297 10608
rect 1177 10536 1221 10570
rect 1255 10536 1297 10570
rect 1177 10498 1297 10536
rect 1177 10464 1221 10498
rect 1255 10464 1297 10498
rect 1177 10426 1297 10464
rect 1177 10392 1221 10426
rect 1255 10392 1297 10426
rect 1177 10334 1297 10392
rect 3916 10766 5155 10810
rect 3916 10334 3964 10766
rect 1177 10290 3964 10334
rect 5104 10334 5155 10766
rect 9753 10748 10992 10800
rect 9753 10334 9802 10748
rect 5104 10290 9802 10334
rect 10942 10334 10992 10748
rect 13697 10790 13817 10828
rect 13697 10756 13739 10790
rect 13773 10756 13817 10790
rect 13697 10718 13817 10756
rect 13697 10684 13739 10718
rect 13773 10684 13817 10718
rect 13697 10646 13817 10684
rect 13697 10612 13739 10646
rect 13773 10612 13817 10646
rect 13697 10574 13817 10612
rect 13697 10540 13739 10574
rect 13773 10540 13817 10574
rect 13697 10502 13817 10540
rect 13697 10468 13739 10502
rect 13773 10468 13817 10502
rect 13697 10430 13817 10468
rect 13697 10396 13739 10430
rect 13773 10396 13817 10430
rect 13697 10334 13817 10396
rect 10942 10290 13817 10334
rect 1177 10256 1355 10290
rect 1389 10256 1427 10290
rect 1461 10256 1499 10290
rect 1533 10256 1571 10290
rect 1605 10256 1643 10290
rect 1677 10256 1715 10290
rect 1749 10256 1787 10290
rect 1821 10256 1859 10290
rect 1893 10256 1931 10290
rect 1965 10256 2003 10290
rect 2037 10256 2075 10290
rect 2109 10256 2147 10290
rect 2181 10256 2219 10290
rect 2253 10256 2291 10290
rect 2325 10256 2363 10290
rect 2397 10256 2435 10290
rect 2469 10256 2507 10290
rect 2541 10256 2579 10290
rect 2613 10256 2651 10290
rect 2685 10256 2723 10290
rect 2757 10256 2795 10290
rect 2829 10256 2867 10290
rect 2901 10256 2939 10290
rect 2973 10256 3011 10290
rect 3045 10256 3083 10290
rect 3117 10256 3155 10290
rect 3189 10256 3227 10290
rect 3261 10256 3299 10290
rect 3333 10256 3371 10290
rect 3405 10256 3443 10290
rect 3477 10256 3515 10290
rect 3549 10256 3587 10290
rect 3621 10256 3659 10290
rect 3693 10256 3731 10290
rect 3765 10256 3803 10290
rect 3837 10256 3875 10290
rect 3909 10256 3947 10290
rect 3981 10256 4019 10266
rect 4053 10256 4091 10266
rect 4125 10256 4163 10266
rect 4197 10256 4235 10266
rect 4269 10256 4307 10266
rect 4341 10256 4379 10266
rect 4413 10256 4451 10266
rect 4485 10256 4523 10266
rect 4557 10256 4595 10266
rect 4629 10256 4667 10266
rect 4701 10256 4739 10266
rect 4773 10256 4811 10266
rect 4845 10256 4883 10266
rect 4917 10256 4955 10266
rect 4989 10256 5027 10266
rect 5061 10256 5099 10266
rect 5133 10256 5171 10290
rect 5205 10256 5243 10290
rect 5277 10256 5315 10290
rect 5349 10256 5387 10290
rect 5421 10256 5459 10290
rect 5493 10256 5531 10290
rect 5565 10256 5603 10290
rect 5637 10256 5675 10290
rect 5709 10256 5747 10290
rect 5781 10256 5819 10290
rect 5853 10256 5891 10290
rect 5925 10256 5963 10290
rect 5997 10256 6035 10290
rect 6069 10256 6107 10290
rect 6141 10256 6179 10290
rect 6213 10256 6251 10290
rect 6285 10256 6323 10290
rect 6357 10256 6395 10290
rect 6429 10256 6467 10290
rect 6501 10256 6539 10290
rect 6573 10256 6611 10290
rect 6645 10256 6683 10290
rect 6717 10256 6755 10290
rect 6789 10256 6827 10290
rect 6861 10256 6899 10290
rect 6933 10256 6971 10290
rect 7005 10256 7043 10290
rect 7077 10256 7115 10290
rect 7149 10256 7187 10290
rect 7221 10256 7259 10290
rect 7293 10256 7331 10290
rect 7365 10256 7403 10290
rect 7437 10256 7475 10290
rect 7509 10256 7547 10290
rect 7581 10256 7619 10290
rect 7653 10256 7691 10290
rect 7725 10256 7763 10290
rect 7797 10256 7835 10290
rect 7869 10256 7907 10290
rect 7941 10256 7979 10290
rect 8013 10256 8051 10290
rect 8085 10256 8123 10290
rect 8157 10256 8195 10290
rect 8229 10256 8267 10290
rect 8301 10256 8339 10290
rect 8373 10256 8411 10290
rect 8445 10256 8483 10290
rect 8517 10256 8555 10290
rect 8589 10256 8627 10290
rect 8661 10256 8699 10290
rect 8733 10256 8771 10290
rect 8805 10256 8843 10290
rect 8877 10256 8915 10290
rect 8949 10256 8987 10290
rect 9021 10256 9059 10290
rect 9093 10256 9131 10290
rect 9165 10256 9203 10290
rect 9237 10256 9275 10290
rect 9309 10256 9347 10290
rect 9381 10256 9419 10290
rect 9453 10256 9491 10290
rect 9525 10256 9563 10290
rect 9597 10256 9635 10290
rect 9669 10256 9707 10290
rect 9741 10256 9779 10290
rect 10965 10256 11003 10290
rect 11037 10256 11075 10290
rect 11109 10256 11147 10290
rect 11181 10256 11219 10290
rect 11253 10256 11291 10290
rect 11325 10256 11363 10290
rect 11397 10256 11435 10290
rect 11469 10256 11507 10290
rect 11541 10256 11579 10290
rect 11613 10256 11651 10290
rect 11685 10256 11723 10290
rect 11757 10256 11795 10290
rect 11829 10256 11867 10290
rect 11901 10256 11939 10290
rect 11973 10256 12011 10290
rect 12045 10256 12083 10290
rect 12117 10256 12155 10290
rect 12189 10256 12227 10290
rect 12261 10256 12299 10290
rect 12333 10256 12371 10290
rect 12405 10256 12443 10290
rect 12477 10256 12515 10290
rect 12549 10256 12587 10290
rect 12621 10256 12659 10290
rect 12693 10256 12731 10290
rect 12765 10256 12803 10290
rect 12837 10256 12875 10290
rect 12909 10256 12947 10290
rect 12981 10256 13019 10290
rect 13053 10256 13091 10290
rect 13125 10256 13163 10290
rect 13197 10256 13235 10290
rect 13269 10256 13307 10290
rect 13341 10256 13379 10290
rect 13413 10256 13451 10290
rect 13485 10256 13523 10290
rect 13557 10256 13595 10290
rect 13629 10256 13817 10290
rect 1177 10248 9802 10256
rect 10942 10248 13817 10256
rect 1177 10214 13817 10248
rect 14099 34680 14219 34718
rect 14099 34646 14120 34680
rect 14154 34646 14219 34680
rect 14099 34608 14219 34646
rect 14099 34574 14120 34608
rect 14154 34574 14219 34608
rect 14099 34536 14219 34574
rect 14099 34502 14120 34536
rect 14154 34502 14219 34536
rect 14099 34464 14219 34502
rect 14099 34430 14120 34464
rect 14154 34430 14219 34464
rect 14099 34392 14219 34430
rect 14099 34358 14120 34392
rect 14154 34358 14219 34392
rect 14099 34320 14219 34358
rect 14099 34286 14120 34320
rect 14154 34286 14219 34320
rect 14099 34248 14219 34286
rect 14099 34214 14120 34248
rect 14154 34214 14219 34248
rect 14099 34176 14219 34214
rect 14099 34142 14120 34176
rect 14154 34142 14219 34176
rect 14099 34104 14219 34142
rect 14099 34070 14120 34104
rect 14154 34070 14219 34104
rect 14099 34032 14219 34070
rect 14099 33998 14120 34032
rect 14154 33998 14219 34032
rect 14099 33960 14219 33998
rect 14099 33926 14120 33960
rect 14154 33926 14219 33960
rect 14099 33888 14219 33926
rect 14099 33854 14120 33888
rect 14154 33854 14219 33888
rect 14099 33816 14219 33854
rect 14099 33782 14120 33816
rect 14154 33782 14219 33816
rect 14099 33744 14219 33782
rect 14099 33710 14120 33744
rect 14154 33710 14219 33744
rect 14099 33672 14219 33710
rect 14099 33638 14120 33672
rect 14154 33638 14219 33672
rect 14099 33600 14219 33638
rect 14099 33566 14120 33600
rect 14154 33566 14219 33600
rect 14099 33528 14219 33566
rect 14099 33494 14120 33528
rect 14154 33494 14219 33528
rect 14099 33456 14219 33494
rect 14099 33422 14120 33456
rect 14154 33422 14219 33456
rect 14099 33384 14219 33422
rect 14099 33350 14120 33384
rect 14154 33350 14219 33384
rect 14099 33312 14219 33350
rect 14099 33278 14120 33312
rect 14154 33278 14219 33312
rect 14099 33240 14219 33278
rect 14099 33206 14120 33240
rect 14154 33206 14219 33240
rect 14099 33168 14219 33206
rect 14099 33134 14120 33168
rect 14154 33134 14219 33168
rect 14099 33096 14219 33134
rect 14099 33062 14120 33096
rect 14154 33062 14219 33096
rect 14099 33024 14219 33062
rect 14099 32990 14120 33024
rect 14154 32990 14219 33024
rect 14099 32952 14219 32990
rect 14099 32918 14120 32952
rect 14154 32918 14219 32952
rect 14099 32880 14219 32918
rect 14099 32846 14120 32880
rect 14154 32846 14219 32880
rect 14099 32808 14219 32846
rect 14099 32774 14120 32808
rect 14154 32774 14219 32808
rect 14099 32736 14219 32774
rect 14099 32702 14120 32736
rect 14154 32702 14219 32736
rect 14099 32664 14219 32702
rect 14099 32630 14120 32664
rect 14154 32630 14219 32664
rect 14099 32592 14219 32630
rect 14099 32558 14120 32592
rect 14154 32558 14219 32592
rect 14099 32520 14219 32558
rect 14099 32486 14120 32520
rect 14154 32486 14219 32520
rect 14099 32448 14219 32486
rect 14099 32414 14120 32448
rect 14154 32414 14219 32448
rect 14099 32376 14219 32414
rect 14099 32342 14120 32376
rect 14154 32342 14219 32376
rect 14099 32304 14219 32342
rect 14099 32270 14120 32304
rect 14154 32270 14219 32304
rect 14099 32232 14219 32270
rect 14099 32198 14120 32232
rect 14154 32198 14219 32232
rect 14099 32160 14219 32198
rect 14099 32126 14120 32160
rect 14154 32126 14219 32160
rect 14099 32088 14219 32126
rect 14099 32054 14120 32088
rect 14154 32054 14219 32088
rect 14099 32016 14219 32054
rect 14099 31982 14120 32016
rect 14154 31982 14219 32016
rect 14099 31944 14219 31982
rect 14099 31910 14120 31944
rect 14154 31910 14219 31944
rect 14099 31872 14219 31910
rect 14099 31838 14120 31872
rect 14154 31838 14219 31872
rect 14099 31800 14219 31838
rect 14099 31766 14120 31800
rect 14154 31766 14219 31800
rect 14099 31728 14219 31766
rect 14099 31694 14120 31728
rect 14154 31694 14219 31728
rect 14099 31656 14219 31694
rect 14099 31622 14120 31656
rect 14154 31622 14219 31656
rect 14099 31584 14219 31622
rect 14099 31550 14120 31584
rect 14154 31550 14219 31584
rect 14099 31512 14219 31550
rect 14099 31478 14120 31512
rect 14154 31478 14219 31512
rect 14099 31440 14219 31478
rect 14099 31406 14120 31440
rect 14154 31406 14219 31440
rect 14099 31368 14219 31406
rect 14099 31334 14120 31368
rect 14154 31334 14219 31368
rect 14099 31296 14219 31334
rect 14099 31262 14120 31296
rect 14154 31262 14219 31296
rect 14099 31224 14219 31262
rect 14099 31190 14120 31224
rect 14154 31190 14219 31224
rect 14099 31152 14219 31190
rect 14099 31118 14120 31152
rect 14154 31118 14219 31152
rect 14099 31080 14219 31118
rect 14099 31046 14120 31080
rect 14154 31046 14219 31080
rect 14099 31008 14219 31046
rect 14099 30974 14120 31008
rect 14154 30974 14219 31008
rect 14099 30936 14219 30974
rect 14099 30902 14120 30936
rect 14154 30902 14219 30936
rect 14099 30864 14219 30902
rect 14099 30830 14120 30864
rect 14154 30830 14219 30864
rect 14099 30792 14219 30830
rect 14099 30758 14120 30792
rect 14154 30758 14219 30792
rect 14099 30720 14219 30758
rect 14099 30686 14120 30720
rect 14154 30686 14219 30720
rect 14099 30648 14219 30686
rect 14099 30614 14120 30648
rect 14154 30614 14219 30648
rect 14099 30576 14219 30614
rect 14099 30542 14120 30576
rect 14154 30542 14219 30576
rect 14099 30504 14219 30542
rect 14099 30470 14120 30504
rect 14154 30470 14219 30504
rect 14099 30432 14219 30470
rect 14099 30398 14120 30432
rect 14154 30398 14219 30432
rect 14099 30360 14219 30398
rect 14099 30326 14120 30360
rect 14154 30326 14219 30360
rect 14099 30288 14219 30326
rect 14099 30254 14120 30288
rect 14154 30254 14219 30288
rect 14099 30216 14219 30254
rect 14099 30182 14120 30216
rect 14154 30182 14219 30216
rect 14099 30144 14219 30182
rect 14099 30110 14120 30144
rect 14154 30110 14219 30144
rect 14099 30072 14219 30110
rect 14099 30038 14120 30072
rect 14154 30038 14219 30072
rect 14099 30000 14219 30038
rect 14099 29966 14120 30000
rect 14154 29966 14219 30000
rect 14099 29928 14219 29966
rect 14099 29894 14120 29928
rect 14154 29894 14219 29928
rect 14099 29856 14219 29894
rect 14099 29822 14120 29856
rect 14154 29822 14219 29856
rect 14099 29784 14219 29822
rect 14099 29750 14120 29784
rect 14154 29750 14219 29784
rect 14099 29712 14219 29750
rect 14099 29678 14120 29712
rect 14154 29678 14219 29712
rect 14099 29640 14219 29678
rect 14099 29606 14120 29640
rect 14154 29606 14219 29640
rect 14099 29568 14219 29606
rect 14099 29534 14120 29568
rect 14154 29534 14219 29568
rect 14099 29496 14219 29534
rect 14099 29462 14120 29496
rect 14154 29462 14219 29496
rect 14099 29424 14219 29462
rect 14099 29390 14120 29424
rect 14154 29390 14219 29424
rect 14099 29352 14219 29390
rect 14099 29318 14120 29352
rect 14154 29318 14219 29352
rect 14099 29280 14219 29318
rect 14099 29246 14120 29280
rect 14154 29246 14219 29280
rect 14099 29208 14219 29246
rect 14099 29174 14120 29208
rect 14154 29174 14219 29208
rect 14099 29136 14219 29174
rect 14099 29102 14120 29136
rect 14154 29102 14219 29136
rect 14099 29064 14219 29102
rect 14099 29030 14120 29064
rect 14154 29030 14219 29064
rect 14099 28992 14219 29030
rect 14099 28958 14120 28992
rect 14154 28958 14219 28992
rect 14099 28920 14219 28958
rect 14099 28886 14120 28920
rect 14154 28886 14219 28920
rect 14099 28848 14219 28886
rect 14099 28814 14120 28848
rect 14154 28814 14219 28848
rect 14099 28776 14219 28814
rect 14099 28742 14120 28776
rect 14154 28742 14219 28776
rect 14099 28704 14219 28742
rect 14099 28670 14120 28704
rect 14154 28670 14219 28704
rect 14099 28632 14219 28670
rect 14099 28598 14120 28632
rect 14154 28598 14219 28632
rect 14099 28560 14219 28598
rect 14099 28526 14120 28560
rect 14154 28526 14219 28560
rect 14099 28488 14219 28526
rect 14099 28454 14120 28488
rect 14154 28454 14219 28488
rect 14099 28416 14219 28454
rect 14099 28382 14120 28416
rect 14154 28382 14219 28416
rect 14099 28344 14219 28382
rect 14099 28310 14120 28344
rect 14154 28310 14219 28344
rect 14099 28272 14219 28310
rect 14099 28238 14120 28272
rect 14154 28238 14219 28272
rect 14099 28200 14219 28238
rect 14099 28166 14120 28200
rect 14154 28166 14219 28200
rect 14099 28128 14219 28166
rect 14099 28094 14120 28128
rect 14154 28094 14219 28128
rect 14099 28056 14219 28094
rect 14099 28022 14120 28056
rect 14154 28022 14219 28056
rect 14099 27984 14219 28022
rect 14099 27950 14120 27984
rect 14154 27950 14219 27984
rect 14099 27912 14219 27950
rect 14099 27878 14120 27912
rect 14154 27878 14219 27912
rect 14099 27840 14219 27878
rect 14099 27806 14120 27840
rect 14154 27806 14219 27840
rect 14099 27768 14219 27806
rect 14099 27734 14120 27768
rect 14154 27734 14219 27768
rect 14099 27696 14219 27734
rect 14099 27662 14120 27696
rect 14154 27662 14219 27696
rect 14099 27624 14219 27662
rect 14099 27590 14120 27624
rect 14154 27590 14219 27624
rect 14099 27552 14219 27590
rect 14099 27518 14120 27552
rect 14154 27518 14219 27552
rect 14099 27480 14219 27518
rect 14099 27446 14120 27480
rect 14154 27446 14219 27480
rect 14099 27408 14219 27446
rect 14099 27374 14120 27408
rect 14154 27374 14219 27408
rect 14099 27336 14219 27374
rect 14099 27302 14120 27336
rect 14154 27302 14219 27336
rect 14099 27264 14219 27302
rect 14099 27230 14120 27264
rect 14154 27230 14219 27264
rect 14099 27192 14219 27230
rect 14099 27158 14120 27192
rect 14154 27158 14219 27192
rect 14099 27120 14219 27158
rect 14099 27086 14120 27120
rect 14154 27086 14219 27120
rect 14099 27048 14219 27086
rect 14099 27014 14120 27048
rect 14154 27014 14219 27048
rect 14099 26976 14219 27014
rect 14099 26942 14120 26976
rect 14154 26942 14219 26976
rect 14099 26904 14219 26942
rect 14099 26870 14120 26904
rect 14154 26870 14219 26904
rect 14099 26832 14219 26870
rect 14099 26798 14120 26832
rect 14154 26798 14219 26832
rect 14099 26760 14219 26798
rect 14099 26726 14120 26760
rect 14154 26726 14219 26760
rect 14099 26688 14219 26726
rect 14099 26654 14120 26688
rect 14154 26654 14219 26688
rect 14099 26616 14219 26654
rect 14099 26582 14120 26616
rect 14154 26582 14219 26616
rect 14099 26544 14219 26582
rect 14099 26510 14120 26544
rect 14154 26510 14219 26544
rect 14099 26472 14219 26510
rect 14099 26438 14120 26472
rect 14154 26438 14219 26472
rect 14099 26400 14219 26438
rect 14099 26366 14120 26400
rect 14154 26366 14219 26400
rect 14099 26328 14219 26366
rect 14099 26294 14120 26328
rect 14154 26294 14219 26328
rect 14099 26256 14219 26294
rect 14099 26222 14120 26256
rect 14154 26222 14219 26256
rect 14099 26184 14219 26222
rect 14099 26150 14120 26184
rect 14154 26150 14219 26184
rect 14099 26112 14219 26150
rect 14099 26078 14120 26112
rect 14154 26078 14219 26112
rect 14099 26040 14219 26078
rect 14099 26006 14120 26040
rect 14154 26006 14219 26040
rect 14099 25968 14219 26006
rect 14099 25934 14120 25968
rect 14154 25934 14219 25968
rect 14099 25896 14219 25934
rect 14099 25862 14120 25896
rect 14154 25862 14219 25896
rect 14099 25824 14219 25862
rect 14099 25790 14120 25824
rect 14154 25790 14219 25824
rect 14099 25752 14219 25790
rect 14099 25718 14120 25752
rect 14154 25718 14219 25752
rect 14099 25680 14219 25718
rect 14099 25646 14120 25680
rect 14154 25646 14219 25680
rect 14099 25608 14219 25646
rect 14099 25574 14120 25608
rect 14154 25574 14219 25608
rect 14099 25536 14219 25574
rect 14099 25502 14120 25536
rect 14154 25502 14219 25536
rect 14099 25464 14219 25502
rect 14099 25430 14120 25464
rect 14154 25430 14219 25464
rect 14099 25392 14219 25430
rect 14099 25358 14120 25392
rect 14154 25358 14219 25392
rect 14099 25320 14219 25358
rect 14099 25286 14120 25320
rect 14154 25286 14219 25320
rect 14099 25248 14219 25286
rect 14099 25214 14120 25248
rect 14154 25214 14219 25248
rect 14099 25176 14219 25214
rect 14099 25142 14120 25176
rect 14154 25142 14219 25176
rect 14099 25104 14219 25142
rect 14099 25070 14120 25104
rect 14154 25070 14219 25104
rect 14099 25032 14219 25070
rect 14099 24998 14120 25032
rect 14154 24998 14219 25032
rect 14099 24960 14219 24998
rect 14099 24926 14120 24960
rect 14154 24926 14219 24960
rect 14099 24888 14219 24926
rect 14099 24854 14120 24888
rect 14154 24854 14219 24888
rect 14099 24816 14219 24854
rect 14099 24782 14120 24816
rect 14154 24782 14219 24816
rect 14099 24744 14219 24782
rect 14099 24710 14120 24744
rect 14154 24710 14219 24744
rect 14099 24672 14219 24710
rect 14099 24638 14120 24672
rect 14154 24638 14219 24672
rect 14099 24600 14219 24638
rect 14099 24566 14120 24600
rect 14154 24566 14219 24600
rect 14099 24528 14219 24566
rect 14099 24494 14120 24528
rect 14154 24494 14219 24528
rect 14099 24456 14219 24494
rect 14099 24422 14120 24456
rect 14154 24422 14219 24456
rect 14099 24384 14219 24422
rect 14099 24350 14120 24384
rect 14154 24350 14219 24384
rect 14099 24312 14219 24350
rect 14099 24278 14120 24312
rect 14154 24278 14219 24312
rect 14099 24240 14219 24278
rect 14099 24206 14120 24240
rect 14154 24206 14219 24240
rect 14099 24168 14219 24206
rect 14099 24134 14120 24168
rect 14154 24134 14219 24168
rect 14099 24096 14219 24134
rect 14099 24062 14120 24096
rect 14154 24062 14219 24096
rect 14099 24024 14219 24062
rect 14099 23990 14120 24024
rect 14154 23990 14219 24024
rect 14099 23952 14219 23990
rect 14099 23918 14120 23952
rect 14154 23918 14219 23952
rect 14099 23880 14219 23918
rect 14099 23846 14120 23880
rect 14154 23846 14219 23880
rect 14099 23808 14219 23846
rect 14099 23774 14120 23808
rect 14154 23774 14219 23808
rect 14099 23736 14219 23774
rect 14099 23702 14120 23736
rect 14154 23702 14219 23736
rect 14099 23664 14219 23702
rect 14099 23630 14120 23664
rect 14154 23630 14219 23664
rect 14099 23592 14219 23630
rect 14099 23558 14120 23592
rect 14154 23558 14219 23592
rect 14099 23520 14219 23558
rect 14099 23486 14120 23520
rect 14154 23486 14219 23520
rect 14099 23448 14219 23486
rect 14099 23414 14120 23448
rect 14154 23414 14219 23448
rect 14099 23376 14219 23414
rect 14099 23342 14120 23376
rect 14154 23342 14219 23376
rect 14099 23304 14219 23342
rect 14099 23270 14120 23304
rect 14154 23270 14219 23304
rect 14099 23232 14219 23270
rect 14099 23198 14120 23232
rect 14154 23198 14219 23232
rect 14099 23160 14219 23198
rect 14099 23126 14120 23160
rect 14154 23126 14219 23160
rect 14099 23088 14219 23126
rect 14099 23054 14120 23088
rect 14154 23054 14219 23088
rect 14099 23016 14219 23054
rect 14099 22982 14120 23016
rect 14154 22982 14219 23016
rect 14099 22944 14219 22982
rect 14099 22910 14120 22944
rect 14154 22910 14219 22944
rect 14099 22872 14219 22910
rect 14099 22838 14120 22872
rect 14154 22838 14219 22872
rect 14099 22800 14219 22838
rect 14099 22766 14120 22800
rect 14154 22766 14219 22800
rect 14099 22728 14219 22766
rect 14099 22694 14120 22728
rect 14154 22694 14219 22728
rect 14099 22656 14219 22694
rect 14099 22622 14120 22656
rect 14154 22622 14219 22656
rect 14099 22584 14219 22622
rect 14099 22550 14120 22584
rect 14154 22550 14219 22584
rect 14099 22512 14219 22550
rect 14099 22478 14120 22512
rect 14154 22478 14219 22512
rect 14099 22440 14219 22478
rect 14099 22406 14120 22440
rect 14154 22406 14219 22440
rect 14099 22368 14219 22406
rect 14099 22334 14120 22368
rect 14154 22334 14219 22368
rect 14099 22296 14219 22334
rect 14099 22262 14120 22296
rect 14154 22262 14219 22296
rect 14099 22224 14219 22262
rect 14099 22190 14120 22224
rect 14154 22190 14219 22224
rect 14099 22152 14219 22190
rect 14099 22118 14120 22152
rect 14154 22118 14219 22152
rect 14099 22080 14219 22118
rect 14099 22046 14120 22080
rect 14154 22046 14219 22080
rect 14099 22008 14219 22046
rect 14099 21974 14120 22008
rect 14154 21974 14219 22008
rect 14099 21936 14219 21974
rect 14099 21902 14120 21936
rect 14154 21902 14219 21936
rect 14099 21864 14219 21902
rect 14099 21830 14120 21864
rect 14154 21830 14219 21864
rect 14099 21792 14219 21830
rect 14099 21758 14120 21792
rect 14154 21758 14219 21792
rect 14099 21720 14219 21758
rect 14099 21686 14120 21720
rect 14154 21686 14219 21720
rect 14099 21648 14219 21686
rect 14099 21614 14120 21648
rect 14154 21614 14219 21648
rect 14099 21576 14219 21614
rect 14099 21542 14120 21576
rect 14154 21542 14219 21576
rect 14099 21504 14219 21542
rect 14099 21470 14120 21504
rect 14154 21470 14219 21504
rect 14099 21432 14219 21470
rect 14099 21398 14120 21432
rect 14154 21398 14219 21432
rect 14099 21360 14219 21398
rect 14099 21326 14120 21360
rect 14154 21326 14219 21360
rect 14099 21288 14219 21326
rect 14099 21254 14120 21288
rect 14154 21254 14219 21288
rect 14099 21216 14219 21254
rect 14099 21182 14120 21216
rect 14154 21182 14219 21216
rect 14099 21144 14219 21182
rect 14099 21110 14120 21144
rect 14154 21110 14219 21144
rect 14099 21072 14219 21110
rect 14099 21038 14120 21072
rect 14154 21038 14219 21072
rect 14099 21000 14219 21038
rect 14099 20966 14120 21000
rect 14154 20966 14219 21000
rect 14099 20928 14219 20966
rect 14099 20894 14120 20928
rect 14154 20894 14219 20928
rect 14099 20856 14219 20894
rect 14099 20822 14120 20856
rect 14154 20822 14219 20856
rect 14099 20784 14219 20822
rect 14099 20750 14120 20784
rect 14154 20750 14219 20784
rect 14099 20712 14219 20750
rect 14099 20678 14120 20712
rect 14154 20678 14219 20712
rect 14099 20640 14219 20678
rect 14099 20606 14120 20640
rect 14154 20606 14219 20640
rect 14099 20568 14219 20606
rect 14099 20534 14120 20568
rect 14154 20534 14219 20568
rect 14099 20496 14219 20534
rect 14099 20462 14120 20496
rect 14154 20462 14219 20496
rect 14099 20424 14219 20462
rect 14099 20390 14120 20424
rect 14154 20390 14219 20424
rect 14099 20352 14219 20390
rect 14099 20318 14120 20352
rect 14154 20318 14219 20352
rect 14099 20280 14219 20318
rect 14099 20246 14120 20280
rect 14154 20246 14219 20280
rect 14099 20208 14219 20246
rect 14099 20174 14120 20208
rect 14154 20174 14219 20208
rect 14099 20136 14219 20174
rect 14099 20102 14120 20136
rect 14154 20102 14219 20136
rect 14099 20064 14219 20102
rect 14099 20030 14120 20064
rect 14154 20030 14219 20064
rect 14099 19992 14219 20030
rect 14099 19958 14120 19992
rect 14154 19958 14219 19992
rect 14099 19920 14219 19958
rect 14099 19886 14120 19920
rect 14154 19886 14219 19920
rect 14099 19848 14219 19886
rect 14099 19814 14120 19848
rect 14154 19814 14219 19848
rect 14099 19776 14219 19814
rect 14099 19742 14120 19776
rect 14154 19742 14219 19776
rect 14099 19704 14219 19742
rect 14099 19670 14120 19704
rect 14154 19670 14219 19704
rect 14099 19632 14219 19670
rect 14099 19598 14120 19632
rect 14154 19598 14219 19632
rect 14099 19560 14219 19598
rect 14099 19526 14120 19560
rect 14154 19526 14219 19560
rect 14099 19488 14219 19526
rect 14099 19454 14120 19488
rect 14154 19454 14219 19488
rect 14099 19416 14219 19454
rect 14099 19382 14120 19416
rect 14154 19382 14219 19416
rect 14099 19344 14219 19382
rect 14099 19310 14120 19344
rect 14154 19310 14219 19344
rect 14099 19272 14219 19310
rect 14099 19238 14120 19272
rect 14154 19238 14219 19272
rect 14099 19200 14219 19238
rect 14099 19166 14120 19200
rect 14154 19166 14219 19200
rect 14099 19128 14219 19166
rect 14099 19094 14120 19128
rect 14154 19094 14219 19128
rect 14099 19056 14219 19094
rect 14099 19022 14120 19056
rect 14154 19022 14219 19056
rect 14099 18984 14219 19022
rect 14099 18950 14120 18984
rect 14154 18950 14219 18984
rect 14099 18912 14219 18950
rect 14099 18878 14120 18912
rect 14154 18878 14219 18912
rect 14099 18840 14219 18878
rect 14099 18806 14120 18840
rect 14154 18806 14219 18840
rect 14099 18768 14219 18806
rect 14099 18734 14120 18768
rect 14154 18734 14219 18768
rect 14099 18696 14219 18734
rect 14099 18662 14120 18696
rect 14154 18662 14219 18696
rect 14099 18624 14219 18662
rect 14099 18590 14120 18624
rect 14154 18590 14219 18624
rect 14099 18552 14219 18590
rect 14099 18518 14120 18552
rect 14154 18518 14219 18552
rect 14099 18480 14219 18518
rect 14099 18446 14120 18480
rect 14154 18446 14219 18480
rect 14099 18408 14219 18446
rect 14099 18374 14120 18408
rect 14154 18374 14219 18408
rect 14099 18336 14219 18374
rect 14099 18302 14120 18336
rect 14154 18302 14219 18336
rect 14099 18264 14219 18302
rect 14099 18230 14120 18264
rect 14154 18230 14219 18264
rect 14099 18192 14219 18230
rect 14099 18158 14120 18192
rect 14154 18158 14219 18192
rect 14099 18120 14219 18158
rect 14099 18086 14120 18120
rect 14154 18086 14219 18120
rect 14099 18048 14219 18086
rect 14099 18014 14120 18048
rect 14154 18014 14219 18048
rect 14099 17976 14219 18014
rect 14099 17942 14120 17976
rect 14154 17942 14219 17976
rect 14099 17904 14219 17942
rect 14099 17870 14120 17904
rect 14154 17870 14219 17904
rect 14099 17832 14219 17870
rect 14099 17798 14120 17832
rect 14154 17798 14219 17832
rect 14099 17760 14219 17798
rect 14099 17726 14120 17760
rect 14154 17726 14219 17760
rect 14099 17688 14219 17726
rect 14099 17654 14120 17688
rect 14154 17654 14219 17688
rect 14099 17616 14219 17654
rect 14099 17582 14120 17616
rect 14154 17582 14219 17616
rect 14099 17544 14219 17582
rect 14099 17510 14120 17544
rect 14154 17510 14219 17544
rect 14099 17472 14219 17510
rect 14099 17438 14120 17472
rect 14154 17438 14219 17472
rect 14099 17400 14219 17438
rect 14099 17366 14120 17400
rect 14154 17366 14219 17400
rect 14099 17328 14219 17366
rect 14099 17294 14120 17328
rect 14154 17294 14219 17328
rect 14099 17256 14219 17294
rect 14099 17222 14120 17256
rect 14154 17222 14219 17256
rect 14099 17184 14219 17222
rect 14099 17150 14120 17184
rect 14154 17150 14219 17184
rect 14099 17112 14219 17150
rect 14099 17078 14120 17112
rect 14154 17078 14219 17112
rect 14099 17040 14219 17078
rect 14099 17006 14120 17040
rect 14154 17006 14219 17040
rect 14099 16968 14219 17006
rect 14099 16934 14120 16968
rect 14154 16934 14219 16968
rect 14099 16896 14219 16934
rect 14099 16862 14120 16896
rect 14154 16862 14219 16896
rect 14099 16824 14219 16862
rect 14099 16790 14120 16824
rect 14154 16790 14219 16824
rect 14099 16752 14219 16790
rect 14099 16718 14120 16752
rect 14154 16718 14219 16752
rect 14099 16680 14219 16718
rect 14099 16646 14120 16680
rect 14154 16646 14219 16680
rect 14099 16608 14219 16646
rect 14099 16574 14120 16608
rect 14154 16574 14219 16608
rect 14099 16536 14219 16574
rect 14099 16502 14120 16536
rect 14154 16502 14219 16536
rect 14099 16464 14219 16502
rect 14099 16430 14120 16464
rect 14154 16430 14219 16464
rect 14099 16392 14219 16430
rect 14099 16358 14120 16392
rect 14154 16358 14219 16392
rect 14099 16320 14219 16358
rect 14099 16286 14120 16320
rect 14154 16286 14219 16320
rect 14099 16248 14219 16286
rect 14099 16214 14120 16248
rect 14154 16214 14219 16248
rect 14099 16176 14219 16214
rect 14099 16142 14120 16176
rect 14154 16142 14219 16176
rect 14099 16104 14219 16142
rect 14099 16070 14120 16104
rect 14154 16070 14219 16104
rect 14099 16032 14219 16070
rect 14099 15998 14120 16032
rect 14154 15998 14219 16032
rect 14099 15960 14219 15998
rect 14099 15926 14120 15960
rect 14154 15926 14219 15960
rect 14099 15888 14219 15926
rect 14099 15854 14120 15888
rect 14154 15854 14219 15888
rect 14099 15816 14219 15854
rect 14099 15782 14120 15816
rect 14154 15782 14219 15816
rect 14099 15744 14219 15782
rect 14099 15710 14120 15744
rect 14154 15710 14219 15744
rect 14099 15672 14219 15710
rect 14099 15638 14120 15672
rect 14154 15638 14219 15672
rect 14099 15600 14219 15638
rect 14099 15566 14120 15600
rect 14154 15566 14219 15600
rect 14099 15528 14219 15566
rect 14099 15494 14120 15528
rect 14154 15494 14219 15528
rect 14099 15456 14219 15494
rect 14099 15422 14120 15456
rect 14154 15422 14219 15456
rect 14099 15384 14219 15422
rect 14099 15350 14120 15384
rect 14154 15350 14219 15384
rect 14099 15312 14219 15350
rect 14099 15278 14120 15312
rect 14154 15278 14219 15312
rect 14099 15240 14219 15278
rect 14099 15206 14120 15240
rect 14154 15206 14219 15240
rect 14099 15168 14219 15206
rect 14099 15134 14120 15168
rect 14154 15134 14219 15168
rect 14099 15096 14219 15134
rect 14099 15062 14120 15096
rect 14154 15062 14219 15096
rect 14099 15024 14219 15062
rect 14099 14990 14120 15024
rect 14154 14990 14219 15024
rect 14099 14952 14219 14990
rect 14099 14918 14120 14952
rect 14154 14918 14219 14952
rect 14099 14880 14219 14918
rect 14099 14846 14120 14880
rect 14154 14846 14219 14880
rect 14099 14808 14219 14846
rect 14099 14774 14120 14808
rect 14154 14774 14219 14808
rect 14099 14736 14219 14774
rect 14099 14702 14120 14736
rect 14154 14702 14219 14736
rect 14099 14664 14219 14702
rect 14099 14630 14120 14664
rect 14154 14630 14219 14664
rect 14099 14592 14219 14630
rect 14099 14558 14120 14592
rect 14154 14558 14219 14592
rect 14099 14520 14219 14558
rect 14099 14486 14120 14520
rect 14154 14486 14219 14520
rect 14099 14448 14219 14486
rect 14099 14414 14120 14448
rect 14154 14414 14219 14448
rect 14099 14376 14219 14414
rect 14099 14342 14120 14376
rect 14154 14342 14219 14376
rect 14099 14304 14219 14342
rect 14099 14270 14120 14304
rect 14154 14270 14219 14304
rect 14099 14232 14219 14270
rect 14099 14198 14120 14232
rect 14154 14198 14219 14232
rect 14099 14160 14219 14198
rect 14099 14126 14120 14160
rect 14154 14126 14219 14160
rect 14099 14088 14219 14126
rect 14099 14054 14120 14088
rect 14154 14054 14219 14088
rect 14099 14016 14219 14054
rect 14099 13982 14120 14016
rect 14154 13982 14219 14016
rect 14099 13944 14219 13982
rect 14099 13910 14120 13944
rect 14154 13910 14219 13944
rect 14099 13872 14219 13910
rect 14099 13838 14120 13872
rect 14154 13838 14219 13872
rect 14099 13800 14219 13838
rect 14099 13766 14120 13800
rect 14154 13766 14219 13800
rect 14099 13728 14219 13766
rect 14099 13694 14120 13728
rect 14154 13694 14219 13728
rect 14099 13656 14219 13694
rect 14099 13622 14120 13656
rect 14154 13622 14219 13656
rect 14099 13584 14219 13622
rect 14099 13550 14120 13584
rect 14154 13550 14219 13584
rect 14099 13512 14219 13550
rect 14099 13478 14120 13512
rect 14154 13478 14219 13512
rect 14099 13440 14219 13478
rect 14099 13406 14120 13440
rect 14154 13406 14219 13440
rect 14099 13368 14219 13406
rect 14099 13334 14120 13368
rect 14154 13334 14219 13368
rect 14099 13296 14219 13334
rect 14099 13262 14120 13296
rect 14154 13262 14219 13296
rect 14099 13224 14219 13262
rect 14099 13190 14120 13224
rect 14154 13190 14219 13224
rect 14099 13152 14219 13190
rect 14099 13118 14120 13152
rect 14154 13118 14219 13152
rect 14099 13080 14219 13118
rect 14099 13046 14120 13080
rect 14154 13046 14219 13080
rect 14099 13008 14219 13046
rect 14099 12974 14120 13008
rect 14154 12974 14219 13008
rect 14099 12936 14219 12974
rect 14099 12902 14120 12936
rect 14154 12902 14219 12936
rect 14099 12864 14219 12902
rect 14099 12830 14120 12864
rect 14154 12830 14219 12864
rect 14099 12792 14219 12830
rect 14099 12758 14120 12792
rect 14154 12758 14219 12792
rect 14099 12720 14219 12758
rect 14099 12686 14120 12720
rect 14154 12686 14219 12720
rect 14099 12648 14219 12686
rect 14099 12614 14120 12648
rect 14154 12614 14219 12648
rect 14099 12576 14219 12614
rect 14099 12542 14120 12576
rect 14154 12542 14219 12576
rect 14099 12504 14219 12542
rect 14099 12470 14120 12504
rect 14154 12470 14219 12504
rect 14099 12432 14219 12470
rect 14099 12398 14120 12432
rect 14154 12398 14219 12432
rect 14099 12360 14219 12398
rect 14099 12326 14120 12360
rect 14154 12326 14219 12360
rect 14099 12288 14219 12326
rect 14099 12254 14120 12288
rect 14154 12254 14219 12288
rect 14099 12216 14219 12254
rect 14099 12182 14120 12216
rect 14154 12182 14219 12216
rect 14099 12144 14219 12182
rect 14099 12110 14120 12144
rect 14154 12110 14219 12144
rect 14099 12072 14219 12110
rect 14099 12038 14120 12072
rect 14154 12038 14219 12072
rect 14099 12000 14219 12038
rect 14099 11966 14120 12000
rect 14154 11966 14219 12000
rect 14099 11928 14219 11966
rect 14099 11894 14120 11928
rect 14154 11894 14219 11928
rect 14099 11856 14219 11894
rect 14099 11822 14120 11856
rect 14154 11822 14219 11856
rect 14099 11784 14219 11822
rect 14099 11750 14120 11784
rect 14154 11750 14219 11784
rect 14099 11712 14219 11750
rect 14099 11678 14120 11712
rect 14154 11678 14219 11712
rect 14099 11640 14219 11678
rect 14099 11606 14120 11640
rect 14154 11606 14219 11640
rect 14099 11568 14219 11606
rect 14099 11534 14120 11568
rect 14154 11534 14219 11568
rect 14099 11496 14219 11534
rect 14099 11462 14120 11496
rect 14154 11462 14219 11496
rect 14099 11424 14219 11462
rect 14099 11390 14120 11424
rect 14154 11390 14219 11424
rect 14099 11352 14219 11390
rect 14099 11318 14120 11352
rect 14154 11318 14219 11352
rect 14099 11280 14219 11318
rect 14099 11246 14120 11280
rect 14154 11246 14219 11280
rect 14099 11208 14219 11246
rect 14099 11174 14120 11208
rect 14154 11174 14219 11208
rect 14099 11136 14219 11174
rect 14099 11102 14120 11136
rect 14154 11102 14219 11136
rect 14099 11064 14219 11102
rect 14099 11030 14120 11064
rect 14154 11030 14219 11064
rect 14099 10992 14219 11030
rect 14099 10958 14120 10992
rect 14154 10958 14219 10992
rect 14099 10920 14219 10958
rect 14099 10886 14120 10920
rect 14154 10886 14219 10920
rect 14099 10848 14219 10886
rect 14099 10814 14120 10848
rect 14154 10814 14219 10848
rect 14099 10776 14219 10814
rect 14099 10742 14120 10776
rect 14154 10742 14219 10776
rect 14099 10704 14219 10742
rect 14099 10670 14120 10704
rect 14154 10670 14219 10704
rect 14099 10632 14219 10670
rect 14099 10598 14120 10632
rect 14154 10598 14219 10632
rect 14099 10560 14219 10598
rect 14099 10526 14120 10560
rect 14154 10526 14219 10560
rect 14099 10488 14219 10526
rect 14099 10454 14120 10488
rect 14154 10454 14219 10488
rect 14099 10416 14219 10454
rect 14099 10382 14120 10416
rect 14154 10382 14219 10416
rect 14099 10344 14219 10382
rect 14099 10310 14120 10344
rect 14154 10310 14219 10344
rect 14099 10272 14219 10310
rect 14099 10238 14120 10272
rect 14154 10238 14219 10272
rect 9753 10209 10992 10214
rect 757 10173 814 10207
rect 848 10173 877 10207
rect 757 10135 877 10173
rect 757 10101 814 10135
rect 848 10101 877 10135
rect 757 9982 877 10101
rect 14099 10200 14219 10238
rect 14099 10166 14120 10200
rect 14154 10166 14219 10200
rect 14099 10128 14219 10166
rect 14099 10094 14120 10128
rect 14154 10094 14219 10128
tri 877 9982 898 10003 sw
tri 14078 9982 14099 10003 se
rect 14099 9982 14219 10094
rect 757 9963 898 9982
tri 898 9963 917 9982 sw
tri 14059 9963 14078 9982 se
rect 14078 9963 14219 9982
rect 757 9943 14219 9963
tri 757 9942 758 9943 ne
rect 758 9942 14186 9943
rect 245 9879 320 9913
rect 354 9879 430 9913
tri 758 9908 792 9942 ne
rect 792 9908 912 9942
rect 946 9908 984 9942
rect 1018 9908 1056 9942
rect 1090 9908 1128 9942
rect 1162 9908 1200 9942
rect 1234 9908 1272 9942
rect 1306 9908 1344 9942
rect 1378 9908 1416 9942
rect 1450 9908 1488 9942
rect 1522 9908 1560 9942
rect 1594 9908 1632 9942
rect 1666 9908 1704 9942
rect 1738 9908 1776 9942
rect 1810 9908 1848 9942
rect 1882 9908 1920 9942
rect 1954 9908 1992 9942
rect 2026 9908 2064 9942
rect 2098 9908 2136 9942
rect 2170 9908 2208 9942
rect 2242 9908 2280 9942
rect 2314 9908 2352 9942
rect 2386 9908 2424 9942
rect 2458 9908 2496 9942
rect 2530 9908 2568 9942
rect 2602 9908 2640 9942
rect 2674 9908 2712 9942
rect 2746 9908 2784 9942
rect 2818 9908 2856 9942
rect 2890 9908 2928 9942
rect 2962 9908 3000 9942
rect 3034 9908 3072 9942
rect 3106 9908 3144 9942
rect 3178 9908 3216 9942
rect 3250 9908 3288 9942
rect 3322 9908 3360 9942
rect 3394 9908 3432 9942
rect 3466 9908 3504 9942
rect 3538 9908 3576 9942
rect 3610 9908 3648 9942
rect 3682 9908 3720 9942
rect 3754 9908 3792 9942
rect 3826 9908 3864 9942
rect 3898 9908 3936 9942
rect 3970 9908 4008 9942
rect 4042 9908 4080 9942
rect 4114 9908 4152 9942
rect 4186 9908 4224 9942
rect 4258 9908 4296 9942
rect 4330 9908 4368 9942
rect 4402 9908 4440 9942
rect 4474 9908 4512 9942
rect 4546 9908 4584 9942
rect 4618 9908 4656 9942
rect 4690 9908 4728 9942
rect 4762 9908 4800 9942
rect 4834 9908 4872 9942
rect 4906 9908 4944 9942
rect 4978 9908 5016 9942
rect 5050 9908 5088 9942
rect 5122 9908 5160 9942
rect 5194 9908 5232 9942
rect 5266 9908 5304 9942
rect 5338 9908 5376 9942
rect 5410 9908 5448 9942
rect 5482 9908 5520 9942
rect 5554 9908 5592 9942
rect 5626 9908 5664 9942
rect 5698 9908 5736 9942
rect 5770 9908 5808 9942
rect 5842 9908 5880 9942
rect 5914 9908 5952 9942
rect 5986 9908 6024 9942
rect 6058 9908 6096 9942
rect 6130 9908 6168 9942
rect 6202 9908 6240 9942
rect 6274 9908 6312 9942
rect 6346 9908 6384 9942
rect 6418 9908 6456 9942
rect 6490 9908 6528 9942
rect 6562 9908 6600 9942
rect 6634 9908 6672 9942
rect 6706 9908 6744 9942
rect 6778 9908 6816 9942
rect 6850 9908 6888 9942
rect 6922 9908 6960 9942
rect 6994 9908 7032 9942
rect 7066 9908 7104 9942
rect 7138 9908 7176 9942
rect 7210 9908 7248 9942
rect 7282 9908 7320 9942
rect 7354 9908 7392 9942
rect 7426 9908 7464 9942
rect 7498 9908 7536 9942
rect 7570 9908 7608 9942
rect 7642 9908 7680 9942
rect 7714 9908 7752 9942
rect 7786 9908 7824 9942
rect 7858 9908 7896 9942
rect 7930 9908 7968 9942
rect 8002 9908 8040 9942
rect 8074 9908 8112 9942
rect 8146 9908 8184 9942
rect 8218 9908 8256 9942
rect 8290 9908 8328 9942
rect 8362 9908 8400 9942
rect 8434 9908 8472 9942
rect 8506 9908 8544 9942
rect 8578 9908 8616 9942
rect 8650 9908 8688 9942
rect 8722 9908 8760 9942
rect 8794 9908 8832 9942
rect 8866 9908 8904 9942
rect 8938 9908 8976 9942
rect 9010 9908 9048 9942
rect 9082 9908 9120 9942
rect 9154 9908 9192 9942
rect 9226 9908 9264 9942
rect 9298 9908 9336 9942
rect 9370 9908 9408 9942
rect 9442 9908 9480 9942
rect 9514 9908 9552 9942
rect 9586 9908 9624 9942
rect 9658 9908 9696 9942
rect 9730 9908 9768 9942
rect 9802 9908 9840 9942
rect 9874 9908 9912 9942
rect 9946 9908 9984 9942
rect 10018 9908 10056 9942
rect 10090 9908 10128 9942
rect 10162 9908 10200 9942
rect 10234 9908 10272 9942
rect 10306 9908 10344 9942
rect 10378 9908 10416 9942
rect 10450 9908 10488 9942
rect 10522 9908 10560 9942
rect 10594 9908 10632 9942
rect 10666 9908 10704 9942
rect 10738 9908 10776 9942
rect 10810 9908 10848 9942
rect 10882 9908 10920 9942
rect 10954 9908 10992 9942
rect 11026 9908 11064 9942
rect 11098 9908 11136 9942
rect 11170 9908 11208 9942
rect 11242 9908 11280 9942
rect 11314 9908 11352 9942
rect 11386 9908 11424 9942
rect 11458 9908 11496 9942
rect 11530 9908 11568 9942
rect 11602 9908 11640 9942
rect 11674 9908 11712 9942
rect 11746 9908 11784 9942
rect 11818 9908 11856 9942
rect 11890 9908 11928 9942
rect 11962 9908 12000 9942
rect 12034 9908 12072 9942
rect 12106 9908 12144 9942
rect 12178 9908 12216 9942
rect 12250 9908 12288 9942
rect 12322 9908 12360 9942
rect 12394 9908 12432 9942
rect 12466 9908 12504 9942
rect 12538 9908 12576 9942
rect 12610 9908 12648 9942
rect 12682 9908 12720 9942
rect 12754 9908 12792 9942
rect 12826 9908 12864 9942
rect 12898 9908 12936 9942
rect 12970 9908 13008 9942
rect 13042 9908 13080 9942
rect 13114 9908 13152 9942
rect 13186 9908 13224 9942
rect 13258 9908 13296 9942
rect 13330 9908 13368 9942
rect 13402 9908 13440 9942
rect 13474 9908 13512 9942
rect 13546 9908 13584 9942
rect 13618 9908 13656 9942
rect 13690 9908 13728 9942
rect 13762 9908 13800 9942
rect 13834 9908 13872 9942
rect 13906 9908 13944 9942
rect 13978 9908 14016 9942
rect 14050 9910 14186 9942
tri 14186 9910 14219 9943 nw
rect 14539 35940 14614 35974
rect 14648 35940 14724 35974
rect 14539 35902 14724 35940
rect 14539 35868 14614 35902
rect 14648 35868 14724 35902
rect 14539 35830 14724 35868
rect 14539 35796 14614 35830
rect 14648 35796 14724 35830
rect 14539 35758 14724 35796
rect 14539 35724 14614 35758
rect 14648 35724 14724 35758
rect 14539 35686 14724 35724
rect 14539 35652 14614 35686
rect 14648 35652 14724 35686
rect 14539 35614 14724 35652
rect 14539 35580 14614 35614
rect 14648 35580 14724 35614
rect 14539 35542 14724 35580
rect 14539 35508 14614 35542
rect 14648 35508 14724 35542
rect 14539 35470 14724 35508
rect 14539 35436 14614 35470
rect 14648 35436 14724 35470
rect 14539 35398 14724 35436
rect 14539 35364 14614 35398
rect 14648 35364 14724 35398
rect 14539 35326 14724 35364
rect 14539 35292 14614 35326
rect 14648 35292 14724 35326
rect 14539 35254 14724 35292
rect 14539 35220 14614 35254
rect 14648 35220 14724 35254
rect 14539 35182 14724 35220
rect 14539 35148 14614 35182
rect 14648 35148 14724 35182
rect 14539 35110 14724 35148
rect 14539 35076 14614 35110
rect 14648 35076 14724 35110
rect 14539 35038 14724 35076
rect 14539 35004 14614 35038
rect 14648 35004 14724 35038
rect 14539 34966 14724 35004
rect 14539 34932 14614 34966
rect 14648 34932 14724 34966
rect 14539 34894 14724 34932
rect 14539 34860 14614 34894
rect 14648 34860 14724 34894
rect 14539 34822 14724 34860
rect 14539 34788 14614 34822
rect 14648 34788 14724 34822
rect 14539 34750 14724 34788
rect 14539 34716 14614 34750
rect 14648 34716 14724 34750
rect 14539 34678 14724 34716
rect 14539 34644 14614 34678
rect 14648 34644 14724 34678
rect 14539 34606 14724 34644
rect 14539 34572 14614 34606
rect 14648 34572 14724 34606
rect 14539 34534 14724 34572
rect 14539 34500 14614 34534
rect 14648 34500 14724 34534
rect 14539 34462 14724 34500
rect 14539 34428 14614 34462
rect 14648 34428 14724 34462
rect 14539 34390 14724 34428
rect 14539 34356 14614 34390
rect 14648 34356 14724 34390
rect 14539 34318 14724 34356
rect 14539 34284 14614 34318
rect 14648 34284 14724 34318
rect 14539 34246 14724 34284
rect 14539 34212 14614 34246
rect 14648 34212 14724 34246
rect 14539 34174 14724 34212
rect 14539 34140 14614 34174
rect 14648 34140 14724 34174
rect 14539 34102 14724 34140
rect 14539 34068 14614 34102
rect 14648 34068 14724 34102
rect 14539 34030 14724 34068
rect 14539 33996 14614 34030
rect 14648 33996 14724 34030
rect 14539 33958 14724 33996
rect 14539 33924 14614 33958
rect 14648 33924 14724 33958
rect 14539 33886 14724 33924
rect 14539 33852 14614 33886
rect 14648 33852 14724 33886
rect 14539 33814 14724 33852
rect 14539 33780 14614 33814
rect 14648 33780 14724 33814
rect 14539 33742 14724 33780
rect 14539 33708 14614 33742
rect 14648 33708 14724 33742
rect 14539 33670 14724 33708
rect 14539 33636 14614 33670
rect 14648 33636 14724 33670
rect 14539 33598 14724 33636
rect 14539 33564 14614 33598
rect 14648 33564 14724 33598
rect 14539 33526 14724 33564
rect 14539 33492 14614 33526
rect 14648 33492 14724 33526
rect 14539 33454 14724 33492
rect 14539 33420 14614 33454
rect 14648 33420 14724 33454
rect 14539 33382 14724 33420
rect 14539 33348 14614 33382
rect 14648 33348 14724 33382
rect 14539 33310 14724 33348
rect 14539 33276 14614 33310
rect 14648 33276 14724 33310
rect 14539 33238 14724 33276
rect 14539 33204 14614 33238
rect 14648 33204 14724 33238
rect 14539 33166 14724 33204
rect 14539 33132 14614 33166
rect 14648 33132 14724 33166
rect 14539 33094 14724 33132
rect 14539 33060 14614 33094
rect 14648 33060 14724 33094
rect 14539 33022 14724 33060
rect 14539 32988 14614 33022
rect 14648 32988 14724 33022
rect 14539 32950 14724 32988
rect 14539 32916 14614 32950
rect 14648 32916 14724 32950
rect 14539 32878 14724 32916
rect 14539 32844 14614 32878
rect 14648 32844 14724 32878
rect 14539 32806 14724 32844
rect 14539 32772 14614 32806
rect 14648 32772 14724 32806
rect 14539 32734 14724 32772
rect 14539 32700 14614 32734
rect 14648 32700 14724 32734
rect 14539 32662 14724 32700
rect 14539 32628 14614 32662
rect 14648 32628 14724 32662
rect 14539 32590 14724 32628
rect 14539 32556 14614 32590
rect 14648 32556 14724 32590
rect 14539 32518 14724 32556
rect 14539 32484 14614 32518
rect 14648 32484 14724 32518
rect 14539 32446 14724 32484
rect 14539 32412 14614 32446
rect 14648 32412 14724 32446
rect 14539 32374 14724 32412
rect 14539 32340 14614 32374
rect 14648 32340 14724 32374
rect 14539 32302 14724 32340
rect 14539 32268 14614 32302
rect 14648 32268 14724 32302
rect 14539 32230 14724 32268
rect 14539 32196 14614 32230
rect 14648 32196 14724 32230
rect 14539 32158 14724 32196
rect 14539 32124 14614 32158
rect 14648 32124 14724 32158
rect 14539 32086 14724 32124
rect 14539 32052 14614 32086
rect 14648 32052 14724 32086
rect 14539 32014 14724 32052
rect 14539 31980 14614 32014
rect 14648 31980 14724 32014
rect 14539 31942 14724 31980
rect 14539 31908 14614 31942
rect 14648 31908 14724 31942
rect 14539 31870 14724 31908
rect 14539 31836 14614 31870
rect 14648 31836 14724 31870
rect 14539 31798 14724 31836
rect 14539 31764 14614 31798
rect 14648 31764 14724 31798
rect 14539 31726 14724 31764
rect 14539 31692 14614 31726
rect 14648 31692 14724 31726
rect 14539 31654 14724 31692
rect 14539 31620 14614 31654
rect 14648 31620 14724 31654
rect 14539 31582 14724 31620
rect 14539 31548 14614 31582
rect 14648 31548 14724 31582
rect 14539 31510 14724 31548
rect 14539 31476 14614 31510
rect 14648 31476 14724 31510
rect 14539 31438 14724 31476
rect 14539 31404 14614 31438
rect 14648 31404 14724 31438
rect 14539 31366 14724 31404
rect 14539 31332 14614 31366
rect 14648 31332 14724 31366
rect 14539 31294 14724 31332
rect 14539 31260 14614 31294
rect 14648 31260 14724 31294
rect 14539 31222 14724 31260
rect 14539 31188 14614 31222
rect 14648 31188 14724 31222
rect 14539 31150 14724 31188
rect 14539 31116 14614 31150
rect 14648 31116 14724 31150
rect 14539 31078 14724 31116
rect 14539 31044 14614 31078
rect 14648 31044 14724 31078
rect 14539 31006 14724 31044
rect 14539 30972 14614 31006
rect 14648 30972 14724 31006
rect 14539 30934 14724 30972
rect 14539 30900 14614 30934
rect 14648 30900 14724 30934
rect 14539 30862 14724 30900
rect 14539 30828 14614 30862
rect 14648 30828 14724 30862
rect 14539 30790 14724 30828
rect 14539 30756 14614 30790
rect 14648 30756 14724 30790
rect 14539 30718 14724 30756
rect 14539 30684 14614 30718
rect 14648 30684 14724 30718
rect 14539 30646 14724 30684
rect 14539 30612 14614 30646
rect 14648 30612 14724 30646
rect 14539 30574 14724 30612
rect 14539 30540 14614 30574
rect 14648 30540 14724 30574
rect 14539 30502 14724 30540
rect 14539 30468 14614 30502
rect 14648 30468 14724 30502
rect 14539 30430 14724 30468
rect 14539 30396 14614 30430
rect 14648 30396 14724 30430
rect 14539 30358 14724 30396
rect 14539 30324 14614 30358
rect 14648 30324 14724 30358
rect 14539 30286 14724 30324
rect 14539 30252 14614 30286
rect 14648 30252 14724 30286
rect 14539 30214 14724 30252
rect 14539 30180 14614 30214
rect 14648 30180 14724 30214
rect 14539 30142 14724 30180
rect 14539 30108 14614 30142
rect 14648 30108 14724 30142
rect 14539 30070 14724 30108
rect 14539 30036 14614 30070
rect 14648 30036 14724 30070
rect 14539 29998 14724 30036
rect 14539 29964 14614 29998
rect 14648 29964 14724 29998
rect 14539 29926 14724 29964
rect 14539 29892 14614 29926
rect 14648 29892 14724 29926
rect 14539 29854 14724 29892
rect 14539 29820 14614 29854
rect 14648 29820 14724 29854
rect 14539 29782 14724 29820
rect 14539 29748 14614 29782
rect 14648 29748 14724 29782
rect 14539 29710 14724 29748
rect 14539 29676 14614 29710
rect 14648 29676 14724 29710
rect 14539 29638 14724 29676
rect 14539 29604 14614 29638
rect 14648 29604 14724 29638
rect 14539 29566 14724 29604
rect 14539 29532 14614 29566
rect 14648 29532 14724 29566
rect 14539 29494 14724 29532
rect 14539 29460 14614 29494
rect 14648 29460 14724 29494
rect 14539 29422 14724 29460
rect 14539 29388 14614 29422
rect 14648 29388 14724 29422
rect 14539 29350 14724 29388
rect 14539 29316 14614 29350
rect 14648 29316 14724 29350
rect 14539 29278 14724 29316
rect 14539 29244 14614 29278
rect 14648 29244 14724 29278
rect 14539 29206 14724 29244
rect 14539 29172 14614 29206
rect 14648 29172 14724 29206
rect 14539 29134 14724 29172
rect 14539 29100 14614 29134
rect 14648 29100 14724 29134
rect 14539 29062 14724 29100
rect 14539 29028 14614 29062
rect 14648 29028 14724 29062
rect 14539 28990 14724 29028
rect 14539 28956 14614 28990
rect 14648 28956 14724 28990
rect 14539 28918 14724 28956
rect 14539 28884 14614 28918
rect 14648 28884 14724 28918
rect 14539 28846 14724 28884
rect 14539 28812 14614 28846
rect 14648 28812 14724 28846
rect 14539 28774 14724 28812
rect 14539 28740 14614 28774
rect 14648 28740 14724 28774
rect 14539 28702 14724 28740
rect 14539 28668 14614 28702
rect 14648 28668 14724 28702
rect 14539 28630 14724 28668
rect 14539 28596 14614 28630
rect 14648 28596 14724 28630
rect 14539 28558 14724 28596
rect 14539 28524 14614 28558
rect 14648 28524 14724 28558
rect 14539 28486 14724 28524
rect 14539 28452 14614 28486
rect 14648 28452 14724 28486
rect 14539 28414 14724 28452
rect 14539 28380 14614 28414
rect 14648 28380 14724 28414
rect 14539 28342 14724 28380
rect 14539 28308 14614 28342
rect 14648 28308 14724 28342
rect 14539 28270 14724 28308
rect 14539 28236 14614 28270
rect 14648 28236 14724 28270
rect 14539 28198 14724 28236
rect 14539 28164 14614 28198
rect 14648 28164 14724 28198
rect 14539 28126 14724 28164
rect 14539 28092 14614 28126
rect 14648 28092 14724 28126
rect 14539 28054 14724 28092
rect 14539 28020 14614 28054
rect 14648 28020 14724 28054
rect 14539 27982 14724 28020
rect 14539 27948 14614 27982
rect 14648 27948 14724 27982
rect 14539 27910 14724 27948
rect 14539 27876 14614 27910
rect 14648 27876 14724 27910
rect 14539 27838 14724 27876
rect 14539 27804 14614 27838
rect 14648 27804 14724 27838
rect 14539 27766 14724 27804
rect 14539 27732 14614 27766
rect 14648 27732 14724 27766
rect 14539 27694 14724 27732
rect 14539 27660 14614 27694
rect 14648 27660 14724 27694
rect 14539 27622 14724 27660
rect 14539 27588 14614 27622
rect 14648 27588 14724 27622
rect 14539 27550 14724 27588
rect 14539 27516 14614 27550
rect 14648 27516 14724 27550
rect 14539 27478 14724 27516
rect 14539 27444 14614 27478
rect 14648 27444 14724 27478
rect 14539 27406 14724 27444
rect 14539 27372 14614 27406
rect 14648 27372 14724 27406
rect 14539 27334 14724 27372
rect 14539 27300 14614 27334
rect 14648 27300 14724 27334
rect 14539 27262 14724 27300
rect 14539 27228 14614 27262
rect 14648 27228 14724 27262
rect 14539 27190 14724 27228
rect 14539 27156 14614 27190
rect 14648 27156 14724 27190
rect 14539 27118 14724 27156
rect 14539 27084 14614 27118
rect 14648 27084 14724 27118
rect 14539 27046 14724 27084
rect 14539 27012 14614 27046
rect 14648 27012 14724 27046
rect 14539 26974 14724 27012
rect 14539 26940 14614 26974
rect 14648 26940 14724 26974
rect 14539 26902 14724 26940
rect 14539 26868 14614 26902
rect 14648 26868 14724 26902
rect 14539 26830 14724 26868
rect 14539 26796 14614 26830
rect 14648 26796 14724 26830
rect 14539 26758 14724 26796
rect 14539 26724 14614 26758
rect 14648 26724 14724 26758
rect 14539 26686 14724 26724
rect 14539 26652 14614 26686
rect 14648 26652 14724 26686
rect 14539 26614 14724 26652
rect 14539 26580 14614 26614
rect 14648 26580 14724 26614
rect 14539 26542 14724 26580
rect 14539 26508 14614 26542
rect 14648 26508 14724 26542
rect 14539 26470 14724 26508
rect 14539 26436 14614 26470
rect 14648 26436 14724 26470
rect 14539 26398 14724 26436
rect 14539 26364 14614 26398
rect 14648 26364 14724 26398
rect 14539 26326 14724 26364
rect 14539 26292 14614 26326
rect 14648 26292 14724 26326
rect 14539 26254 14724 26292
rect 14539 26220 14614 26254
rect 14648 26220 14724 26254
rect 14539 26182 14724 26220
rect 14539 26148 14614 26182
rect 14648 26148 14724 26182
rect 14539 26110 14724 26148
rect 14539 26076 14614 26110
rect 14648 26076 14724 26110
rect 14539 26038 14724 26076
rect 14539 26004 14614 26038
rect 14648 26004 14724 26038
rect 14539 25966 14724 26004
rect 14539 25932 14614 25966
rect 14648 25932 14724 25966
rect 14539 25894 14724 25932
rect 14539 25860 14614 25894
rect 14648 25860 14724 25894
rect 14539 25822 14724 25860
rect 14539 25788 14614 25822
rect 14648 25788 14724 25822
rect 14539 25750 14724 25788
rect 14539 25716 14614 25750
rect 14648 25716 14724 25750
rect 14539 25678 14724 25716
rect 14539 25644 14614 25678
rect 14648 25644 14724 25678
rect 14539 25606 14724 25644
rect 14539 25572 14614 25606
rect 14648 25572 14724 25606
rect 14539 25534 14724 25572
rect 14539 25500 14614 25534
rect 14648 25500 14724 25534
rect 14539 25462 14724 25500
rect 14539 25428 14614 25462
rect 14648 25428 14724 25462
rect 14539 25390 14724 25428
rect 14539 25356 14614 25390
rect 14648 25356 14724 25390
rect 14539 25318 14724 25356
rect 14539 25284 14614 25318
rect 14648 25284 14724 25318
rect 14539 25246 14724 25284
rect 14539 25212 14614 25246
rect 14648 25212 14724 25246
rect 14539 25174 14724 25212
rect 14539 25140 14614 25174
rect 14648 25140 14724 25174
rect 14539 25102 14724 25140
rect 14539 25068 14614 25102
rect 14648 25068 14724 25102
rect 14539 25030 14724 25068
rect 14539 24996 14614 25030
rect 14648 24996 14724 25030
rect 14539 24958 14724 24996
rect 14539 24924 14614 24958
rect 14648 24924 14724 24958
rect 14539 24886 14724 24924
rect 14539 24852 14614 24886
rect 14648 24852 14724 24886
rect 14539 24814 14724 24852
rect 14539 24780 14614 24814
rect 14648 24780 14724 24814
rect 14539 24742 14724 24780
rect 14539 24708 14614 24742
rect 14648 24708 14724 24742
rect 14539 24670 14724 24708
rect 14539 24636 14614 24670
rect 14648 24636 14724 24670
rect 14539 24598 14724 24636
rect 14539 24564 14614 24598
rect 14648 24564 14724 24598
rect 14539 24526 14724 24564
rect 14539 24492 14614 24526
rect 14648 24492 14724 24526
rect 14539 24454 14724 24492
rect 14539 24420 14614 24454
rect 14648 24420 14724 24454
rect 14539 24382 14724 24420
rect 14539 24348 14614 24382
rect 14648 24348 14724 24382
rect 14539 24310 14724 24348
rect 14539 24276 14614 24310
rect 14648 24276 14724 24310
rect 14539 24238 14724 24276
rect 14539 24204 14614 24238
rect 14648 24204 14724 24238
rect 14539 24166 14724 24204
rect 14539 24132 14614 24166
rect 14648 24132 14724 24166
rect 14539 24094 14724 24132
rect 14539 24060 14614 24094
rect 14648 24060 14724 24094
rect 14539 24022 14724 24060
rect 14539 23988 14614 24022
rect 14648 23988 14724 24022
rect 14539 23950 14724 23988
rect 14539 23916 14614 23950
rect 14648 23916 14724 23950
rect 14539 23878 14724 23916
rect 14539 23844 14614 23878
rect 14648 23844 14724 23878
rect 14539 23806 14724 23844
rect 14539 23772 14614 23806
rect 14648 23772 14724 23806
rect 14539 23734 14724 23772
rect 14539 23700 14614 23734
rect 14648 23700 14724 23734
rect 14539 23662 14724 23700
rect 14539 23628 14614 23662
rect 14648 23628 14724 23662
rect 14539 23590 14724 23628
rect 14539 23556 14614 23590
rect 14648 23556 14724 23590
rect 14539 23518 14724 23556
rect 14539 23484 14614 23518
rect 14648 23484 14724 23518
rect 14539 23446 14724 23484
rect 14539 23412 14614 23446
rect 14648 23412 14724 23446
rect 14539 23374 14724 23412
rect 14539 23340 14614 23374
rect 14648 23340 14724 23374
rect 14539 23302 14724 23340
rect 14539 23268 14614 23302
rect 14648 23268 14724 23302
rect 14539 23230 14724 23268
rect 14539 23196 14614 23230
rect 14648 23196 14724 23230
rect 14539 23158 14724 23196
rect 14539 23124 14614 23158
rect 14648 23124 14724 23158
rect 14539 23086 14724 23124
rect 14539 23052 14614 23086
rect 14648 23052 14724 23086
rect 14539 23014 14724 23052
rect 14539 22980 14614 23014
rect 14648 22980 14724 23014
rect 14539 22942 14724 22980
rect 14539 22908 14614 22942
rect 14648 22908 14724 22942
rect 14539 22870 14724 22908
rect 14539 22836 14614 22870
rect 14648 22836 14724 22870
rect 14539 22798 14724 22836
rect 14539 22764 14614 22798
rect 14648 22764 14724 22798
rect 14539 22726 14724 22764
rect 14539 22692 14614 22726
rect 14648 22692 14724 22726
rect 14539 22654 14724 22692
rect 14539 22620 14614 22654
rect 14648 22620 14724 22654
rect 14539 22582 14724 22620
rect 14539 22548 14614 22582
rect 14648 22548 14724 22582
rect 14539 22510 14724 22548
rect 14539 22476 14614 22510
rect 14648 22476 14724 22510
rect 14539 22438 14724 22476
rect 14539 22404 14614 22438
rect 14648 22404 14724 22438
rect 14539 22366 14724 22404
rect 14539 22332 14614 22366
rect 14648 22332 14724 22366
rect 14539 22294 14724 22332
rect 14539 22260 14614 22294
rect 14648 22260 14724 22294
rect 14539 22222 14724 22260
rect 14539 22188 14614 22222
rect 14648 22188 14724 22222
rect 14539 22150 14724 22188
rect 14539 22116 14614 22150
rect 14648 22116 14724 22150
rect 14539 22078 14724 22116
rect 14539 22044 14614 22078
rect 14648 22044 14724 22078
rect 14539 22006 14724 22044
rect 14539 21972 14614 22006
rect 14648 21972 14724 22006
rect 14539 21934 14724 21972
rect 14539 21900 14614 21934
rect 14648 21900 14724 21934
rect 14539 21862 14724 21900
rect 14539 21828 14614 21862
rect 14648 21828 14724 21862
rect 14539 21790 14724 21828
rect 14539 21756 14614 21790
rect 14648 21756 14724 21790
rect 14539 21718 14724 21756
rect 14539 21684 14614 21718
rect 14648 21684 14724 21718
rect 14539 21646 14724 21684
rect 14539 21612 14614 21646
rect 14648 21612 14724 21646
rect 14539 21574 14724 21612
rect 14539 21540 14614 21574
rect 14648 21540 14724 21574
rect 14539 21502 14724 21540
rect 14539 21468 14614 21502
rect 14648 21468 14724 21502
rect 14539 21430 14724 21468
rect 14539 21396 14614 21430
rect 14648 21396 14724 21430
rect 14539 21358 14724 21396
rect 14539 21324 14614 21358
rect 14648 21324 14724 21358
rect 14539 21286 14724 21324
rect 14539 21252 14614 21286
rect 14648 21252 14724 21286
rect 14539 21214 14724 21252
rect 14539 21180 14614 21214
rect 14648 21180 14724 21214
rect 14539 21142 14724 21180
rect 14539 21108 14614 21142
rect 14648 21108 14724 21142
rect 14539 21070 14724 21108
rect 14539 21036 14614 21070
rect 14648 21036 14724 21070
rect 14539 20998 14724 21036
rect 14539 20964 14614 20998
rect 14648 20964 14724 20998
rect 14539 20926 14724 20964
rect 14539 20892 14614 20926
rect 14648 20892 14724 20926
rect 14539 20854 14724 20892
rect 14539 20820 14614 20854
rect 14648 20820 14724 20854
rect 14539 20782 14724 20820
rect 14539 20748 14614 20782
rect 14648 20748 14724 20782
rect 14539 20710 14724 20748
rect 14539 20676 14614 20710
rect 14648 20676 14724 20710
rect 14539 20638 14724 20676
rect 14539 20604 14614 20638
rect 14648 20604 14724 20638
rect 14539 20566 14724 20604
rect 14539 20532 14614 20566
rect 14648 20532 14724 20566
rect 14539 20494 14724 20532
rect 14539 20460 14614 20494
rect 14648 20460 14724 20494
rect 14539 20422 14724 20460
rect 14539 20388 14614 20422
rect 14648 20388 14724 20422
rect 14539 20350 14724 20388
rect 14539 20316 14614 20350
rect 14648 20316 14724 20350
rect 14539 20278 14724 20316
rect 14539 20244 14614 20278
rect 14648 20244 14724 20278
rect 14539 20206 14724 20244
rect 14539 20172 14614 20206
rect 14648 20172 14724 20206
rect 14539 20134 14724 20172
rect 14539 20100 14614 20134
rect 14648 20100 14724 20134
rect 14539 20062 14724 20100
rect 14539 20028 14614 20062
rect 14648 20028 14724 20062
rect 14539 19990 14724 20028
rect 14539 19956 14614 19990
rect 14648 19956 14724 19990
rect 14539 19918 14724 19956
rect 14539 19884 14614 19918
rect 14648 19884 14724 19918
rect 14539 19846 14724 19884
rect 14539 19812 14614 19846
rect 14648 19812 14724 19846
rect 14539 19774 14724 19812
rect 14539 19740 14614 19774
rect 14648 19740 14724 19774
rect 14539 19702 14724 19740
rect 14539 19668 14614 19702
rect 14648 19668 14724 19702
rect 14539 19630 14724 19668
rect 14539 19596 14614 19630
rect 14648 19596 14724 19630
rect 14539 19558 14724 19596
rect 14539 19524 14614 19558
rect 14648 19524 14724 19558
rect 14539 19486 14724 19524
rect 14539 19452 14614 19486
rect 14648 19452 14724 19486
rect 14539 19414 14724 19452
rect 14539 19380 14614 19414
rect 14648 19380 14724 19414
rect 14539 19342 14724 19380
rect 14539 19308 14614 19342
rect 14648 19308 14724 19342
rect 14539 19270 14724 19308
rect 14539 19236 14614 19270
rect 14648 19236 14724 19270
rect 14539 19198 14724 19236
rect 14539 19164 14614 19198
rect 14648 19164 14724 19198
rect 14539 19126 14724 19164
rect 14539 19092 14614 19126
rect 14648 19092 14724 19126
rect 14539 19054 14724 19092
rect 14539 19020 14614 19054
rect 14648 19020 14724 19054
rect 14539 18982 14724 19020
rect 14539 18948 14614 18982
rect 14648 18948 14724 18982
rect 14539 18910 14724 18948
rect 14539 18876 14614 18910
rect 14648 18876 14724 18910
rect 14539 18838 14724 18876
rect 14539 18804 14614 18838
rect 14648 18804 14724 18838
rect 14539 18766 14724 18804
rect 14539 18732 14614 18766
rect 14648 18732 14724 18766
rect 14539 18694 14724 18732
rect 14539 18660 14614 18694
rect 14648 18660 14724 18694
rect 14539 18622 14724 18660
rect 14539 18588 14614 18622
rect 14648 18588 14724 18622
rect 14539 18550 14724 18588
rect 14539 18516 14614 18550
rect 14648 18516 14724 18550
rect 14539 18478 14724 18516
rect 14539 18444 14614 18478
rect 14648 18444 14724 18478
rect 14539 18406 14724 18444
rect 14539 18372 14614 18406
rect 14648 18372 14724 18406
rect 14539 18334 14724 18372
rect 14539 18300 14614 18334
rect 14648 18300 14724 18334
rect 14539 18262 14724 18300
rect 14539 18228 14614 18262
rect 14648 18228 14724 18262
rect 14539 18190 14724 18228
rect 14539 18156 14614 18190
rect 14648 18156 14724 18190
rect 14539 18118 14724 18156
rect 14539 18084 14614 18118
rect 14648 18084 14724 18118
rect 14539 18046 14724 18084
rect 14539 18012 14614 18046
rect 14648 18012 14724 18046
rect 14539 17974 14724 18012
rect 14539 17940 14614 17974
rect 14648 17940 14724 17974
rect 14539 17902 14724 17940
rect 14539 17868 14614 17902
rect 14648 17868 14724 17902
rect 14539 17830 14724 17868
rect 14539 17796 14614 17830
rect 14648 17796 14724 17830
rect 14539 17758 14724 17796
rect 14539 17724 14614 17758
rect 14648 17724 14724 17758
rect 14539 17686 14724 17724
rect 14539 17652 14614 17686
rect 14648 17652 14724 17686
rect 14539 17614 14724 17652
rect 14539 17580 14614 17614
rect 14648 17580 14724 17614
rect 14539 17542 14724 17580
rect 14539 17508 14614 17542
rect 14648 17508 14724 17542
rect 14539 17470 14724 17508
rect 14539 17436 14614 17470
rect 14648 17436 14724 17470
rect 14539 17398 14724 17436
rect 14539 17364 14614 17398
rect 14648 17364 14724 17398
rect 14539 17326 14724 17364
rect 14539 17292 14614 17326
rect 14648 17292 14724 17326
rect 14539 17254 14724 17292
rect 14539 17220 14614 17254
rect 14648 17220 14724 17254
rect 14539 17182 14724 17220
rect 14539 17148 14614 17182
rect 14648 17148 14724 17182
rect 14539 17110 14724 17148
rect 14539 17076 14614 17110
rect 14648 17076 14724 17110
rect 14539 17038 14724 17076
rect 14539 17004 14614 17038
rect 14648 17004 14724 17038
rect 14539 16966 14724 17004
rect 14539 16932 14614 16966
rect 14648 16932 14724 16966
rect 14539 16894 14724 16932
rect 14539 16860 14614 16894
rect 14648 16860 14724 16894
rect 14539 16822 14724 16860
rect 14539 16788 14614 16822
rect 14648 16788 14724 16822
rect 14539 16750 14724 16788
rect 14539 16716 14614 16750
rect 14648 16716 14724 16750
rect 14539 16678 14724 16716
rect 14539 16644 14614 16678
rect 14648 16644 14724 16678
rect 14539 16606 14724 16644
rect 14539 16572 14614 16606
rect 14648 16572 14724 16606
rect 14539 16534 14724 16572
rect 14539 16500 14614 16534
rect 14648 16500 14724 16534
rect 14539 16462 14724 16500
rect 14539 16428 14614 16462
rect 14648 16428 14724 16462
rect 14539 16390 14724 16428
rect 14539 16356 14614 16390
rect 14648 16356 14724 16390
rect 14539 16318 14724 16356
rect 14539 16284 14614 16318
rect 14648 16284 14724 16318
rect 14539 16246 14724 16284
rect 14539 16212 14614 16246
rect 14648 16212 14724 16246
rect 14539 16174 14724 16212
rect 14539 16140 14614 16174
rect 14648 16140 14724 16174
rect 14539 16102 14724 16140
rect 14539 16068 14614 16102
rect 14648 16068 14724 16102
rect 14539 16030 14724 16068
rect 14539 15996 14614 16030
rect 14648 15996 14724 16030
rect 14539 15958 14724 15996
rect 14539 15924 14614 15958
rect 14648 15924 14724 15958
rect 14539 15886 14724 15924
rect 14539 15852 14614 15886
rect 14648 15852 14724 15886
rect 14539 15814 14724 15852
rect 14539 15780 14614 15814
rect 14648 15780 14724 15814
rect 14539 15742 14724 15780
rect 14539 15708 14614 15742
rect 14648 15708 14724 15742
rect 14539 15670 14724 15708
rect 14539 15636 14614 15670
rect 14648 15636 14724 15670
rect 14539 15598 14724 15636
rect 14539 15564 14614 15598
rect 14648 15564 14724 15598
rect 14539 15526 14724 15564
rect 14539 15492 14614 15526
rect 14648 15492 14724 15526
rect 14539 15454 14724 15492
rect 14539 15420 14614 15454
rect 14648 15420 14724 15454
rect 14539 15382 14724 15420
rect 14539 15348 14614 15382
rect 14648 15348 14724 15382
rect 14539 15310 14724 15348
rect 14539 15276 14614 15310
rect 14648 15276 14724 15310
rect 14539 15238 14724 15276
rect 14539 15204 14614 15238
rect 14648 15204 14724 15238
rect 14539 15166 14724 15204
rect 14539 15132 14614 15166
rect 14648 15132 14724 15166
rect 14539 15094 14724 15132
rect 14539 15060 14614 15094
rect 14648 15060 14724 15094
rect 14539 15022 14724 15060
rect 14539 14988 14614 15022
rect 14648 14988 14724 15022
rect 14539 14950 14724 14988
rect 14539 14916 14614 14950
rect 14648 14916 14724 14950
rect 14539 14878 14724 14916
rect 14539 14844 14614 14878
rect 14648 14844 14724 14878
rect 14539 14806 14724 14844
rect 14539 14772 14614 14806
rect 14648 14772 14724 14806
rect 14539 14734 14724 14772
rect 14539 14700 14614 14734
rect 14648 14700 14724 14734
rect 14539 14662 14724 14700
rect 14539 14628 14614 14662
rect 14648 14628 14724 14662
rect 14539 14590 14724 14628
rect 14539 14556 14614 14590
rect 14648 14556 14724 14590
rect 14539 14518 14724 14556
rect 14539 14484 14614 14518
rect 14648 14484 14724 14518
rect 14539 14446 14724 14484
rect 14539 14412 14614 14446
rect 14648 14412 14724 14446
rect 14539 14374 14724 14412
rect 14539 14340 14614 14374
rect 14648 14340 14724 14374
rect 14539 14302 14724 14340
rect 14539 14268 14614 14302
rect 14648 14268 14724 14302
rect 14539 14230 14724 14268
rect 14539 14196 14614 14230
rect 14648 14196 14724 14230
rect 14539 14158 14724 14196
rect 14539 14124 14614 14158
rect 14648 14124 14724 14158
rect 14539 14086 14724 14124
rect 14539 14052 14614 14086
rect 14648 14052 14724 14086
rect 14539 14014 14724 14052
rect 14539 13980 14614 14014
rect 14648 13980 14724 14014
rect 14539 13942 14724 13980
rect 14539 13908 14614 13942
rect 14648 13908 14724 13942
rect 14539 13870 14724 13908
rect 14539 13836 14614 13870
rect 14648 13836 14724 13870
rect 14539 13798 14724 13836
rect 14539 13764 14614 13798
rect 14648 13764 14724 13798
rect 14539 13726 14724 13764
rect 14539 13692 14614 13726
rect 14648 13692 14724 13726
rect 14539 13654 14724 13692
rect 14539 13620 14614 13654
rect 14648 13620 14724 13654
rect 14539 13582 14724 13620
rect 14539 13548 14614 13582
rect 14648 13548 14724 13582
rect 14539 13510 14724 13548
rect 14539 13476 14614 13510
rect 14648 13476 14724 13510
rect 14539 13438 14724 13476
rect 14539 13404 14614 13438
rect 14648 13404 14724 13438
rect 14539 13366 14724 13404
rect 14539 13332 14614 13366
rect 14648 13332 14724 13366
rect 14539 13294 14724 13332
rect 14539 13260 14614 13294
rect 14648 13260 14724 13294
rect 14539 13222 14724 13260
rect 14539 13188 14614 13222
rect 14648 13188 14724 13222
rect 14539 13150 14724 13188
rect 14539 13116 14614 13150
rect 14648 13116 14724 13150
rect 14539 13078 14724 13116
rect 14539 13044 14614 13078
rect 14648 13044 14724 13078
rect 14539 13006 14724 13044
rect 14539 12972 14614 13006
rect 14648 12972 14724 13006
rect 14539 12934 14724 12972
rect 14539 12900 14614 12934
rect 14648 12900 14724 12934
rect 14539 12862 14724 12900
rect 14539 12828 14614 12862
rect 14648 12828 14724 12862
rect 14539 12790 14724 12828
rect 14539 12756 14614 12790
rect 14648 12756 14724 12790
rect 14539 12718 14724 12756
rect 14539 12684 14614 12718
rect 14648 12684 14724 12718
rect 14539 12646 14724 12684
rect 14539 12612 14614 12646
rect 14648 12612 14724 12646
rect 14539 12574 14724 12612
rect 14539 12540 14614 12574
rect 14648 12540 14724 12574
rect 14539 12502 14724 12540
rect 14539 12468 14614 12502
rect 14648 12468 14724 12502
rect 14539 12430 14724 12468
rect 14539 12396 14614 12430
rect 14648 12396 14724 12430
rect 14539 12358 14724 12396
rect 14539 12324 14614 12358
rect 14648 12324 14724 12358
rect 14539 12286 14724 12324
rect 14539 12252 14614 12286
rect 14648 12252 14724 12286
rect 14539 12214 14724 12252
rect 14539 12180 14614 12214
rect 14648 12180 14724 12214
rect 14539 12142 14724 12180
rect 14539 12108 14614 12142
rect 14648 12108 14724 12142
rect 14539 12070 14724 12108
rect 14539 12036 14614 12070
rect 14648 12036 14724 12070
rect 14539 11998 14724 12036
rect 14539 11964 14614 11998
rect 14648 11964 14724 11998
rect 14539 11926 14724 11964
rect 14539 11892 14614 11926
rect 14648 11892 14724 11926
rect 14539 11854 14724 11892
rect 14539 11820 14614 11854
rect 14648 11820 14724 11854
rect 14539 11782 14724 11820
rect 14539 11748 14614 11782
rect 14648 11748 14724 11782
rect 14539 11710 14724 11748
rect 14539 11676 14614 11710
rect 14648 11676 14724 11710
rect 14539 11638 14724 11676
rect 14539 11604 14614 11638
rect 14648 11604 14724 11638
rect 14539 11566 14724 11604
rect 14539 11532 14614 11566
rect 14648 11532 14724 11566
rect 14539 11494 14724 11532
rect 14539 11460 14614 11494
rect 14648 11460 14724 11494
rect 14539 11422 14724 11460
rect 14539 11388 14614 11422
rect 14648 11388 14724 11422
rect 14539 11350 14724 11388
rect 14539 11316 14614 11350
rect 14648 11316 14724 11350
rect 14539 11278 14724 11316
rect 14539 11244 14614 11278
rect 14648 11244 14724 11278
rect 14539 11206 14724 11244
rect 14539 11172 14614 11206
rect 14648 11172 14724 11206
rect 14539 11134 14724 11172
rect 14539 11100 14614 11134
rect 14648 11100 14724 11134
rect 14539 11062 14724 11100
rect 14539 11028 14614 11062
rect 14648 11028 14724 11062
rect 14539 10990 14724 11028
rect 14539 10956 14614 10990
rect 14648 10956 14724 10990
rect 14539 10918 14724 10956
rect 14539 10884 14614 10918
rect 14648 10884 14724 10918
rect 14539 10846 14724 10884
rect 14539 10812 14614 10846
rect 14648 10812 14724 10846
rect 14539 10774 14724 10812
rect 14539 10740 14614 10774
rect 14648 10740 14724 10774
rect 14539 10702 14724 10740
rect 14539 10668 14614 10702
rect 14648 10668 14724 10702
rect 14539 10630 14724 10668
rect 14539 10596 14614 10630
rect 14648 10596 14724 10630
rect 14539 10558 14724 10596
rect 14539 10524 14614 10558
rect 14648 10524 14724 10558
rect 14539 10486 14724 10524
rect 14539 10452 14614 10486
rect 14648 10452 14724 10486
rect 14539 10414 14724 10452
rect 14539 10380 14614 10414
rect 14648 10380 14724 10414
rect 14539 10342 14724 10380
rect 14539 10308 14614 10342
rect 14648 10308 14724 10342
rect 14539 10270 14724 10308
rect 14539 10236 14614 10270
rect 14648 10236 14724 10270
rect 14539 10198 14724 10236
rect 14539 10164 14614 10198
rect 14648 10164 14724 10198
rect 14539 10126 14724 10164
rect 14539 10092 14614 10126
rect 14648 10092 14724 10126
rect 14539 10054 14724 10092
rect 14539 10020 14614 10054
rect 14648 10020 14724 10054
rect 14539 9982 14724 10020
rect 14539 9948 14614 9982
rect 14648 9948 14724 9982
rect 14539 9910 14724 9948
rect 14050 9908 14152 9910
tri 792 9907 793 9908 ne
rect 793 9907 14152 9908
rect 245 9841 430 9879
tri 793 9876 824 9907 ne
rect 824 9876 14152 9907
tri 14152 9876 14186 9910 nw
rect 14539 9876 14614 9910
rect 14648 9876 14724 9910
tri 824 9843 857 9876 ne
rect 857 9843 14119 9876
tri 14119 9843 14152 9876 nw
rect 245 9807 320 9841
rect 354 9807 430 9841
rect 245 9769 430 9807
rect 245 9735 320 9769
rect 354 9735 430 9769
rect 245 9697 430 9735
rect 245 9663 320 9697
rect 354 9663 430 9697
rect 245 9528 430 9663
rect 858 9774 2096 9843
rect 858 9740 883 9774
rect 917 9752 955 9774
rect 989 9752 1027 9774
rect 1061 9752 1099 9774
rect 1133 9752 1171 9774
rect 1205 9752 1243 9774
rect 1277 9752 1315 9774
rect 1349 9752 1387 9774
rect 1421 9752 1459 9774
rect 1493 9752 1531 9774
rect 1565 9752 1603 9774
rect 1637 9752 1675 9774
rect 1709 9752 1747 9774
rect 1781 9752 1819 9774
rect 1853 9752 1891 9774
rect 1925 9752 1963 9774
rect 1997 9752 2035 9774
rect 2069 9740 2096 9774
rect 245 9452 720 9528
rect 245 9418 320 9452
rect 354 9418 610 9452
rect 644 9418 720 9452
rect 245 9343 720 9418
rect 858 9316 908 9740
rect 2048 9316 2096 9740
rect 12858 9774 14096 9843
rect 12858 9740 12883 9774
rect 12917 9752 12955 9774
rect 12989 9752 13027 9774
rect 13061 9752 13099 9774
rect 13133 9752 13171 9774
rect 13205 9752 13243 9774
rect 13277 9752 13315 9774
rect 13349 9752 13387 9774
rect 13421 9752 13459 9774
rect 13493 9752 13531 9774
rect 13565 9752 13603 9774
rect 13637 9752 13675 9774
rect 13709 9752 13747 9774
rect 13781 9752 13819 9774
rect 13853 9752 13891 9774
rect 13925 9752 13963 9774
rect 13997 9752 14035 9774
rect 14069 9740 14096 9774
rect 11273 9528 12512 9529
rect 2248 9484 12705 9528
rect 2248 9483 11322 9484
rect 2248 9452 2445 9483
rect 3585 9452 11322 9483
rect 12462 9452 12705 9484
rect 2248 9418 2311 9452
rect 2345 9418 2383 9452
rect 2417 9418 2445 9452
rect 3585 9418 3607 9452
rect 3641 9418 3679 9452
rect 3713 9418 3751 9452
rect 3785 9418 3823 9452
rect 3857 9418 3895 9452
rect 3929 9418 3967 9452
rect 4001 9418 4039 9452
rect 4073 9418 4111 9452
rect 4145 9418 4183 9452
rect 4217 9418 4255 9452
rect 4289 9418 4327 9452
rect 4361 9418 4399 9452
rect 4433 9418 4471 9452
rect 4505 9418 4543 9452
rect 4577 9418 4615 9452
rect 4649 9418 4687 9452
rect 4721 9418 4759 9452
rect 4793 9418 4831 9452
rect 4865 9418 4903 9452
rect 4937 9418 4975 9452
rect 5009 9418 5047 9452
rect 5081 9418 5119 9452
rect 5153 9418 5191 9452
rect 5225 9418 5263 9452
rect 5297 9418 5335 9452
rect 5369 9418 5407 9452
rect 5441 9418 5479 9452
rect 5513 9418 5551 9452
rect 5585 9418 5623 9452
rect 5657 9418 5695 9452
rect 5729 9418 5767 9452
rect 5801 9418 5839 9452
rect 5873 9418 5911 9452
rect 5945 9418 5983 9452
rect 6017 9418 6055 9452
rect 6089 9418 6127 9452
rect 6161 9418 6199 9452
rect 6233 9418 6271 9452
rect 6305 9418 6343 9452
rect 6377 9418 6415 9452
rect 6449 9418 6487 9452
rect 6521 9418 6559 9452
rect 6593 9418 6631 9452
rect 6665 9418 6703 9452
rect 6737 9418 6775 9452
rect 6809 9418 6847 9452
rect 6881 9418 6919 9452
rect 6953 9418 6991 9452
rect 7025 9418 7063 9452
rect 7097 9418 7135 9452
rect 7169 9418 7207 9452
rect 7241 9418 7279 9452
rect 7313 9418 7351 9452
rect 7385 9418 7423 9452
rect 7457 9418 7495 9452
rect 7529 9418 7567 9452
rect 7601 9418 7639 9452
rect 7673 9418 7711 9452
rect 7745 9418 7783 9452
rect 7817 9418 7855 9452
rect 7889 9418 7927 9452
rect 7961 9418 7999 9452
rect 8033 9418 8071 9452
rect 8105 9418 8143 9452
rect 8177 9418 8215 9452
rect 8249 9418 8287 9452
rect 8321 9418 8359 9452
rect 8393 9418 8431 9452
rect 8465 9418 8503 9452
rect 8537 9418 8575 9452
rect 8609 9418 8647 9452
rect 8681 9418 8719 9452
rect 8753 9418 8791 9452
rect 8825 9418 8863 9452
rect 8897 9418 8935 9452
rect 8969 9418 9007 9452
rect 9041 9418 9079 9452
rect 9113 9418 9151 9452
rect 9185 9418 9223 9452
rect 9257 9418 9295 9452
rect 9329 9418 9367 9452
rect 9401 9418 9439 9452
rect 9473 9418 9511 9452
rect 9545 9418 9583 9452
rect 9617 9418 9655 9452
rect 9689 9418 9727 9452
rect 9761 9418 9799 9452
rect 9833 9418 9871 9452
rect 9905 9418 9943 9452
rect 9977 9418 10015 9452
rect 10049 9418 10087 9452
rect 10121 9418 10159 9452
rect 10193 9418 10231 9452
rect 10265 9418 10303 9452
rect 10337 9418 10375 9452
rect 10409 9418 10447 9452
rect 10481 9418 10519 9452
rect 10553 9418 10591 9452
rect 10625 9418 10663 9452
rect 10697 9418 10735 9452
rect 10769 9418 10807 9452
rect 10841 9418 10879 9452
rect 10913 9418 10951 9452
rect 10985 9418 11023 9452
rect 11057 9418 11095 9452
rect 11129 9418 11167 9452
rect 11201 9418 11239 9452
rect 11273 9418 11311 9452
rect 12462 9418 12463 9452
rect 12497 9418 12535 9452
rect 12569 9418 12607 9452
rect 12641 9418 12705 9452
rect 2248 9343 2445 9418
rect 858 9252 2096 9316
rect 2396 8983 2445 9343
rect 3585 9343 11322 9418
rect 3585 8983 3635 9343
rect 2396 8939 3635 8983
rect 11273 8984 11322 9343
rect 12462 9343 12705 9418
rect 12462 8984 12512 9343
rect 12858 9316 12908 9740
rect 14048 9316 14096 9740
rect 14539 9838 14724 9876
rect 14539 9804 14614 9838
rect 14648 9804 14724 9838
rect 14539 9766 14724 9804
rect 14539 9732 14614 9766
rect 14648 9732 14724 9766
rect 14539 9694 14724 9732
rect 14539 9660 14614 9694
rect 14648 9660 14724 9694
rect 14539 9528 14724 9660
rect 14232 9452 14724 9528
rect 14232 9418 14314 9452
rect 14348 9418 14614 9452
rect 14648 9418 14724 9452
rect 14232 9343 14724 9418
rect 12858 9252 14096 9316
rect 11273 8940 12512 8984
<< via1 >>
rect 3964 10290 5104 10766
rect 9802 10290 10942 10748
rect 3964 10266 3981 10290
rect 3981 10266 4019 10290
rect 4019 10266 4053 10290
rect 4053 10266 4091 10290
rect 4091 10266 4125 10290
rect 4125 10266 4163 10290
rect 4163 10266 4197 10290
rect 4197 10266 4235 10290
rect 4235 10266 4269 10290
rect 4269 10266 4307 10290
rect 4307 10266 4341 10290
rect 4341 10266 4379 10290
rect 4379 10266 4413 10290
rect 4413 10266 4451 10290
rect 4451 10266 4485 10290
rect 4485 10266 4523 10290
rect 4523 10266 4557 10290
rect 4557 10266 4595 10290
rect 4595 10266 4629 10290
rect 4629 10266 4667 10290
rect 4667 10266 4701 10290
rect 4701 10266 4739 10290
rect 4739 10266 4773 10290
rect 4773 10266 4811 10290
rect 4811 10266 4845 10290
rect 4845 10266 4883 10290
rect 4883 10266 4917 10290
rect 4917 10266 4955 10290
rect 4955 10266 4989 10290
rect 4989 10266 5027 10290
rect 5027 10266 5061 10290
rect 5061 10266 5099 10290
rect 5099 10266 5104 10290
rect 9802 10256 9813 10290
rect 9813 10256 9851 10290
rect 9851 10256 9885 10290
rect 9885 10256 9923 10290
rect 9923 10256 9957 10290
rect 9957 10256 9995 10290
rect 9995 10256 10029 10290
rect 10029 10256 10067 10290
rect 10067 10256 10101 10290
rect 10101 10256 10139 10290
rect 10139 10256 10173 10290
rect 10173 10256 10211 10290
rect 10211 10256 10245 10290
rect 10245 10256 10283 10290
rect 10283 10256 10317 10290
rect 10317 10256 10355 10290
rect 10355 10256 10389 10290
rect 10389 10256 10427 10290
rect 10427 10256 10461 10290
rect 10461 10256 10499 10290
rect 10499 10256 10533 10290
rect 10533 10256 10571 10290
rect 10571 10256 10605 10290
rect 10605 10256 10643 10290
rect 10643 10256 10677 10290
rect 10677 10256 10715 10290
rect 10715 10256 10749 10290
rect 10749 10256 10787 10290
rect 10787 10256 10821 10290
rect 10821 10256 10859 10290
rect 10859 10256 10893 10290
rect 10893 10256 10931 10290
rect 10931 10256 10942 10290
rect 9802 10248 10942 10256
rect 908 9740 917 9752
rect 917 9740 955 9752
rect 955 9740 989 9752
rect 989 9740 1027 9752
rect 1027 9740 1061 9752
rect 1061 9740 1099 9752
rect 1099 9740 1133 9752
rect 1133 9740 1171 9752
rect 1171 9740 1205 9752
rect 1205 9740 1243 9752
rect 1243 9740 1277 9752
rect 1277 9740 1315 9752
rect 1315 9740 1349 9752
rect 1349 9740 1387 9752
rect 1387 9740 1421 9752
rect 1421 9740 1459 9752
rect 1459 9740 1493 9752
rect 1493 9740 1531 9752
rect 1531 9740 1565 9752
rect 1565 9740 1603 9752
rect 1603 9740 1637 9752
rect 1637 9740 1675 9752
rect 1675 9740 1709 9752
rect 1709 9740 1747 9752
rect 1747 9740 1781 9752
rect 1781 9740 1819 9752
rect 1819 9740 1853 9752
rect 1853 9740 1891 9752
rect 1891 9740 1925 9752
rect 1925 9740 1963 9752
rect 1963 9740 1997 9752
rect 1997 9740 2035 9752
rect 2035 9740 2048 9752
rect 908 9316 2048 9740
rect 12908 9740 12917 9752
rect 12917 9740 12955 9752
rect 12955 9740 12989 9752
rect 12989 9740 13027 9752
rect 13027 9740 13061 9752
rect 13061 9740 13099 9752
rect 13099 9740 13133 9752
rect 13133 9740 13171 9752
rect 13171 9740 13205 9752
rect 13205 9740 13243 9752
rect 13243 9740 13277 9752
rect 13277 9740 13315 9752
rect 13315 9740 13349 9752
rect 13349 9740 13387 9752
rect 13387 9740 13421 9752
rect 13421 9740 13459 9752
rect 13459 9740 13493 9752
rect 13493 9740 13531 9752
rect 13531 9740 13565 9752
rect 13565 9740 13603 9752
rect 13603 9740 13637 9752
rect 13637 9740 13675 9752
rect 13675 9740 13709 9752
rect 13709 9740 13747 9752
rect 13747 9740 13781 9752
rect 13781 9740 13819 9752
rect 13819 9740 13853 9752
rect 13853 9740 13891 9752
rect 13891 9740 13925 9752
rect 13925 9740 13963 9752
rect 13963 9740 13997 9752
rect 13997 9740 14035 9752
rect 14035 9740 14048 9752
rect 2445 9452 3585 9483
rect 11322 9452 12462 9484
rect 2445 9418 2455 9452
rect 2455 9418 2489 9452
rect 2489 9418 2527 9452
rect 2527 9418 2561 9452
rect 2561 9418 2599 9452
rect 2599 9418 2633 9452
rect 2633 9418 2671 9452
rect 2671 9418 2705 9452
rect 2705 9418 2743 9452
rect 2743 9418 2777 9452
rect 2777 9418 2815 9452
rect 2815 9418 2849 9452
rect 2849 9418 2887 9452
rect 2887 9418 2921 9452
rect 2921 9418 2959 9452
rect 2959 9418 2993 9452
rect 2993 9418 3031 9452
rect 3031 9418 3065 9452
rect 3065 9418 3103 9452
rect 3103 9418 3137 9452
rect 3137 9418 3175 9452
rect 3175 9418 3209 9452
rect 3209 9418 3247 9452
rect 3247 9418 3281 9452
rect 3281 9418 3319 9452
rect 3319 9418 3353 9452
rect 3353 9418 3391 9452
rect 3391 9418 3425 9452
rect 3425 9418 3463 9452
rect 3463 9418 3497 9452
rect 3497 9418 3535 9452
rect 3535 9418 3569 9452
rect 3569 9418 3585 9452
rect 11322 9418 11345 9452
rect 11345 9418 11383 9452
rect 11383 9418 11417 9452
rect 11417 9418 11455 9452
rect 11455 9418 11489 9452
rect 11489 9418 11527 9452
rect 11527 9418 11561 9452
rect 11561 9418 11599 9452
rect 11599 9418 11633 9452
rect 11633 9418 11671 9452
rect 11671 9418 11705 9452
rect 11705 9418 11743 9452
rect 11743 9418 11777 9452
rect 11777 9418 11815 9452
rect 11815 9418 11849 9452
rect 11849 9418 11887 9452
rect 11887 9418 11921 9452
rect 11921 9418 11959 9452
rect 11959 9418 11993 9452
rect 11993 9418 12031 9452
rect 12031 9418 12065 9452
rect 12065 9418 12103 9452
rect 12103 9418 12137 9452
rect 12137 9418 12175 9452
rect 12175 9418 12209 9452
rect 12209 9418 12247 9452
rect 12247 9418 12281 9452
rect 12281 9418 12319 9452
rect 12319 9418 12353 9452
rect 12353 9418 12391 9452
rect 12391 9418 12425 9452
rect 12425 9418 12462 9452
rect 2445 8983 3585 9418
rect 11322 8984 12462 9418
rect 12908 9316 14048 9740
<< metal2 >>
rect 3916 10784 5155 10810
rect 3916 10248 3946 10784
rect 5122 10248 5155 10784
rect 3916 10219 5155 10248
rect 9753 10766 10992 10794
rect 9753 10230 9784 10766
rect 10960 10230 10992 10766
rect 9753 10209 10992 10230
rect 858 9756 2096 9787
rect 858 9300 890 9756
rect 2066 9300 2096 9756
rect 12858 9752 14096 9787
rect 12858 9741 12908 9752
rect 14048 9741 14096 9752
rect 858 9252 2096 9300
rect 2396 9501 3635 9528
rect 2396 8965 2427 9501
rect 3603 8965 3635 9501
rect 2396 8939 3635 8965
rect 11273 9502 12512 9529
rect 11273 8966 11304 9502
rect 12480 8966 12512 9502
rect 12858 9285 12890 9741
rect 14066 9285 14096 9741
rect 12858 9252 14096 9285
rect 11273 8940 12512 8966
<< via2 >>
rect 3946 10766 5122 10784
rect 3946 10266 3964 10766
rect 3964 10266 5104 10766
rect 5104 10266 5122 10766
rect 3946 10248 5122 10266
rect 9784 10748 10960 10766
rect 9784 10248 9802 10748
rect 9802 10248 10942 10748
rect 10942 10248 10960 10748
rect 9784 10230 10960 10248
rect 890 9752 2066 9756
rect 890 9316 908 9752
rect 908 9316 2048 9752
rect 2048 9316 2066 9752
rect 890 9300 2066 9316
rect 2427 9483 3603 9501
rect 2427 8983 2445 9483
rect 2445 8983 3585 9483
rect 3585 8983 3603 9483
rect 2427 8965 3603 8983
rect 11304 9484 12480 9502
rect 11304 8984 11322 9484
rect 11322 8984 12462 9484
rect 12462 8984 12480 9484
rect 11304 8966 12480 8984
rect 12890 9316 12908 9741
rect 12908 9316 14048 9741
rect 14048 9316 14066 9741
rect 12890 9285 14066 9316
<< metal3 >>
tri 99 33575 1155 34631 se
rect 1155 34618 3100 34631
rect 1155 34554 2276 34618
rect 2340 34554 2359 34618
rect 2423 34554 2443 34618
rect 2507 34554 2527 34618
rect 2591 34554 2611 34618
rect 2675 34554 3100 34618
rect 1155 34524 3100 34554
rect 1155 34460 2276 34524
rect 2340 34460 2359 34524
rect 2423 34460 2443 34524
rect 2507 34460 2527 34524
rect 2591 34460 2611 34524
rect 2675 34460 3100 34524
rect 1155 34441 3100 34460
rect 1155 34377 2148 34441
rect 2212 34430 3100 34441
rect 2212 34377 2276 34430
rect 1155 34366 2276 34377
rect 2340 34366 2359 34430
rect 2423 34366 2443 34430
rect 2507 34366 2527 34430
rect 2591 34366 2611 34430
rect 2675 34366 3100 34430
rect 1155 34336 3100 34366
rect 1155 34316 2276 34336
rect 1155 34252 2004 34316
rect 2068 34252 2084 34316
rect 2148 34252 2164 34316
rect 2228 34272 2276 34316
rect 2340 34272 2359 34336
rect 2423 34272 2443 34336
rect 2507 34272 2527 34336
rect 2591 34272 2611 34336
rect 2675 34272 3100 34336
rect 2228 34252 3100 34272
rect 1155 34242 3100 34252
rect 1155 34220 2276 34242
rect 1155 34183 2004 34220
rect 1155 34119 1890 34183
rect 1954 34156 2004 34183
rect 2068 34156 2084 34220
rect 2148 34156 2164 34220
rect 2228 34178 2276 34220
rect 2340 34178 2359 34242
rect 2423 34178 2443 34242
rect 2507 34178 2527 34242
rect 2591 34178 2611 34242
rect 2675 34178 3100 34242
rect 2228 34156 3100 34178
rect 1954 34148 3100 34156
rect 1954 34119 2276 34148
rect 1155 34084 2276 34119
rect 2340 34084 2359 34148
rect 2423 34084 2443 34148
rect 2507 34084 2527 34148
rect 2591 34084 2611 34148
rect 2675 34084 3100 34148
rect 1155 34078 3100 34084
rect 1155 34014 1748 34078
rect 1812 34014 1837 34078
rect 1901 34014 1927 34078
rect 1991 34014 2017 34078
rect 2081 34014 2107 34078
rect 2171 34014 3100 34078
rect 1155 34009 3100 34014
rect 1155 33962 2247 34009
rect 1155 33898 1748 33962
rect 1812 33898 1837 33962
rect 1901 33898 1927 33962
rect 1991 33898 2017 33962
rect 2081 33898 2107 33962
rect 2171 33945 2247 33962
rect 2311 33945 3100 34009
rect 2171 33898 3100 33945
rect 1155 33886 3100 33898
rect 1155 33822 1644 33886
rect 1708 33848 3100 33886
rect 1708 33846 2700 33848
rect 1708 33822 1748 33846
rect 1155 33782 1748 33822
rect 1812 33782 1837 33846
rect 1901 33782 1927 33846
rect 1991 33782 2017 33846
rect 2081 33782 2107 33846
rect 2171 33782 2700 33846
rect 1155 33754 2700 33782
rect 1155 33690 1424 33754
rect 1488 33690 1513 33754
rect 1577 33690 1603 33754
rect 1667 33690 1693 33754
rect 1757 33690 1783 33754
rect 1847 33721 2700 33754
rect 1847 33690 1929 33721
rect 1155 33657 1929 33690
rect 1993 33657 2700 33721
rect 1155 33638 2700 33657
rect 1155 33575 1424 33638
rect 99 33574 1424 33575
rect 1488 33574 1513 33638
rect 1577 33574 1603 33638
rect 1667 33574 1693 33638
rect 1757 33574 1783 33638
rect 1847 33574 2700 33638
rect 99 33558 2700 33574
rect 99 33494 1316 33558
rect 1380 33522 2700 33558
rect 1380 33494 1424 33522
rect 99 33458 1424 33494
rect 1488 33458 1513 33522
rect 1577 33458 1603 33522
rect 1667 33458 1693 33522
rect 1757 33458 1783 33522
rect 1847 33458 2700 33522
rect 99 33434 2700 33458
tri 2700 33448 3100 33848 nw
rect 11900 34618 13835 34631
rect 11900 34554 12341 34618
rect 12405 34554 12425 34618
rect 12489 34554 12509 34618
rect 12573 34554 12593 34618
rect 12657 34554 12677 34618
rect 12741 34554 13835 34618
rect 11900 34524 13835 34554
rect 11900 34460 12341 34524
rect 12405 34460 12425 34524
rect 12489 34460 12509 34524
rect 12573 34460 12593 34524
rect 12657 34460 12677 34524
rect 12741 34460 13835 34524
rect 11900 34441 13835 34460
rect 11900 34430 12804 34441
rect 11900 34366 12341 34430
rect 12405 34366 12425 34430
rect 12489 34366 12509 34430
rect 12573 34366 12593 34430
rect 12657 34366 12677 34430
rect 12741 34377 12804 34430
rect 12868 34377 13835 34441
rect 12741 34366 13835 34377
rect 11900 34336 13835 34366
rect 11900 34272 12341 34336
rect 12405 34272 12425 34336
rect 12489 34272 12509 34336
rect 12573 34272 12593 34336
rect 12657 34272 12677 34336
rect 12741 34316 13835 34336
rect 12741 34272 12788 34316
rect 11900 34252 12788 34272
rect 12852 34252 12868 34316
rect 12932 34252 12948 34316
rect 13012 34252 13835 34316
rect 11900 34242 13835 34252
rect 11900 34178 12341 34242
rect 12405 34178 12425 34242
rect 12489 34178 12509 34242
rect 12573 34178 12593 34242
rect 12657 34178 12677 34242
rect 12741 34220 13835 34242
rect 12741 34178 12788 34220
rect 11900 34156 12788 34178
rect 12852 34156 12868 34220
rect 12932 34156 12948 34220
rect 13012 34183 13835 34220
rect 13012 34156 13062 34183
rect 11900 34148 13062 34156
rect 11900 34084 12341 34148
rect 12405 34084 12425 34148
rect 12489 34084 12509 34148
rect 12573 34084 12593 34148
rect 12657 34084 12677 34148
rect 12741 34119 13062 34148
rect 13126 34119 13835 34183
rect 12741 34084 13835 34119
rect 11900 34078 13835 34084
rect 11900 34014 12845 34078
rect 12909 34014 12935 34078
rect 12999 34014 13025 34078
rect 13089 34014 13115 34078
rect 13179 34014 13204 34078
rect 13268 34014 13835 34078
rect 11900 34009 13835 34014
rect 11900 33945 12705 34009
rect 12769 33962 13835 34009
rect 12769 33945 12845 33962
rect 11900 33898 12845 33945
rect 12909 33898 12935 33962
rect 12999 33898 13025 33962
rect 13089 33898 13115 33962
rect 13179 33898 13204 33962
rect 13268 33898 13835 33962
rect 11900 33886 13835 33898
rect 11900 33848 13308 33886
tri 11900 33448 12300 33848 ne
rect 12300 33846 13308 33848
rect 12300 33782 12845 33846
rect 12909 33782 12935 33846
rect 12999 33782 13025 33846
rect 13089 33782 13115 33846
rect 13179 33782 13204 33846
rect 13268 33822 13308 33846
rect 13372 33822 13835 33886
rect 13268 33782 13835 33822
rect 12300 33754 13835 33782
rect 12300 33721 13169 33754
rect 12300 33657 13023 33721
rect 13087 33690 13169 33721
rect 13233 33690 13259 33754
rect 13323 33690 13349 33754
rect 13413 33690 13439 33754
rect 13503 33690 13528 33754
rect 13592 33690 13835 33754
rect 13087 33657 13835 33690
rect 12300 33638 13835 33657
rect 12300 33574 13169 33638
rect 13233 33574 13259 33638
rect 13323 33574 13349 33638
rect 13413 33574 13439 33638
rect 13503 33574 13528 33638
rect 13592 33608 13835 33638
tri 13835 33608 14858 34631 sw
rect 13592 33574 14858 33608
rect 12300 33558 14858 33574
rect 12300 33522 13636 33558
rect 12300 33458 13169 33522
rect 13233 33458 13259 33522
rect 13323 33458 13349 33522
rect 13413 33458 13439 33522
rect 13503 33458 13528 33522
rect 13592 33494 13636 33522
rect 13700 33494 14858 33558
rect 13592 33458 14858 33494
rect 99 33370 1104 33434
rect 1168 33370 1193 33434
rect 1257 33370 1283 33434
rect 1347 33370 1373 33434
rect 1437 33370 1463 33434
rect 1527 33396 2700 33434
rect 1527 33370 1604 33396
rect 99 33332 1604 33370
rect 1668 33332 2700 33396
rect 99 33318 2700 33332
rect 99 33254 1104 33318
rect 1168 33254 1193 33318
rect 1257 33254 1283 33318
rect 1347 33254 1373 33318
rect 1437 33254 1463 33318
rect 1527 33254 2700 33318
rect 99 33202 2700 33254
rect 99 33138 1104 33202
rect 1168 33138 1193 33202
rect 1257 33138 1283 33202
rect 1347 33138 1373 33202
rect 1437 33138 1463 33202
rect 1527 33138 2700 33202
rect 99 33109 2700 33138
rect 99 33045 982 33109
rect 1046 33045 1072 33109
rect 1136 33045 1162 33109
rect 1226 33045 1252 33109
rect 1316 33045 1342 33109
rect 1406 33045 1432 33109
rect 1496 33045 2700 33109
rect 99 33029 2700 33045
rect 99 32965 982 33029
rect 1046 32965 1072 33029
rect 1136 32965 1162 33029
rect 1226 32965 1252 33029
rect 1316 32965 1342 33029
rect 1406 32965 1432 33029
rect 1496 32965 2700 33029
rect 99 32949 2700 32965
rect 99 32885 982 32949
rect 1046 32885 1072 32949
rect 1136 32885 1162 32949
rect 1226 32885 1252 32949
rect 1316 32885 1342 32949
rect 1406 32885 1432 32949
rect 1496 32885 2700 32949
rect 99 32869 2700 32885
rect 99 32805 982 32869
rect 1046 32805 1072 32869
rect 1136 32805 1162 32869
rect 1226 32805 1252 32869
rect 1316 32805 1342 32869
rect 1406 32805 1432 32869
rect 1496 32805 2700 32869
rect 99 32789 2700 32805
rect 99 32725 982 32789
rect 1046 32725 1072 32789
rect 1136 32725 1162 32789
rect 1226 32725 1252 32789
rect 1316 32725 1342 32789
rect 1406 32725 1432 32789
rect 1496 32725 2700 32789
rect 99 32709 2700 32725
rect 99 32645 982 32709
rect 1046 32645 1072 32709
rect 1136 32645 1162 32709
rect 1226 32645 1252 32709
rect 1316 32645 1342 32709
rect 1406 32645 1432 32709
rect 1496 32645 2700 32709
rect 99 32629 2700 32645
rect 99 32565 982 32629
rect 1046 32565 1072 32629
rect 1136 32565 1162 32629
rect 1226 32565 1252 32629
rect 1316 32565 1342 32629
rect 1406 32565 1432 32629
rect 1496 32565 2700 32629
rect 99 32549 2700 32565
rect 99 32485 982 32549
rect 1046 32485 1072 32549
rect 1136 32485 1162 32549
rect 1226 32485 1252 32549
rect 1316 32485 1342 32549
rect 1406 32485 1432 32549
rect 1496 32485 2700 32549
rect 99 32469 2700 32485
rect 99 32405 982 32469
rect 1046 32405 1072 32469
rect 1136 32405 1162 32469
rect 1226 32405 1252 32469
rect 1316 32405 1342 32469
rect 1406 32405 1432 32469
rect 1496 32405 2700 32469
rect 99 32389 2700 32405
rect 99 32325 982 32389
rect 1046 32325 1072 32389
rect 1136 32325 1162 32389
rect 1226 32325 1252 32389
rect 1316 32325 1342 32389
rect 1406 32325 1432 32389
rect 1496 32325 2700 32389
rect 99 32309 2700 32325
rect 99 32245 982 32309
rect 1046 32245 1072 32309
rect 1136 32245 1162 32309
rect 1226 32245 1252 32309
rect 1316 32245 1342 32309
rect 1406 32245 1432 32309
rect 1496 32245 2700 32309
rect 99 32229 2700 32245
rect 99 32165 982 32229
rect 1046 32165 1072 32229
rect 1136 32165 1162 32229
rect 1226 32165 1252 32229
rect 1316 32165 1342 32229
rect 1406 32165 1432 32229
rect 1496 32165 2700 32229
rect 99 32149 2700 32165
rect 99 32085 982 32149
rect 1046 32085 1072 32149
rect 1136 32085 1162 32149
rect 1226 32085 1252 32149
rect 1316 32085 1342 32149
rect 1406 32085 1432 32149
rect 1496 32085 2700 32149
rect 99 32069 2700 32085
rect 99 32005 982 32069
rect 1046 32005 1072 32069
rect 1136 32005 1162 32069
rect 1226 32005 1252 32069
rect 1316 32005 1342 32069
rect 1406 32005 1432 32069
rect 1496 32005 2700 32069
rect 99 31989 2700 32005
rect 99 31925 982 31989
rect 1046 31925 1072 31989
rect 1136 31925 1162 31989
rect 1226 31925 1252 31989
rect 1316 31925 1342 31989
rect 1406 31925 1432 31989
rect 1496 31925 2700 31989
rect 99 31909 2700 31925
rect 99 31845 982 31909
rect 1046 31845 1072 31909
rect 1136 31845 1162 31909
rect 1226 31845 1252 31909
rect 1316 31845 1342 31909
rect 1406 31845 1432 31909
rect 1496 31845 2700 31909
rect 99 31829 2700 31845
rect 99 31765 982 31829
rect 1046 31765 1072 31829
rect 1136 31765 1162 31829
rect 1226 31765 1252 31829
rect 1316 31765 1342 31829
rect 1406 31765 1432 31829
rect 1496 31765 2700 31829
rect 99 31749 2700 31765
rect 99 31685 982 31749
rect 1046 31685 1072 31749
rect 1136 31685 1162 31749
rect 1226 31685 1252 31749
rect 1316 31685 1342 31749
rect 1406 31685 1432 31749
rect 1496 31685 2700 31749
rect 99 31669 2700 31685
rect 99 31605 982 31669
rect 1046 31605 1072 31669
rect 1136 31605 1162 31669
rect 1226 31605 1252 31669
rect 1316 31605 1342 31669
rect 1406 31605 1432 31669
rect 1496 31605 2700 31669
rect 99 31589 2700 31605
rect 99 31525 982 31589
rect 1046 31525 1072 31589
rect 1136 31525 1162 31589
rect 1226 31525 1252 31589
rect 1316 31525 1342 31589
rect 1406 31525 1432 31589
rect 1496 31525 2700 31589
rect 99 31509 2700 31525
rect 99 31445 982 31509
rect 1046 31445 1072 31509
rect 1136 31445 1162 31509
rect 1226 31445 1252 31509
rect 1316 31445 1342 31509
rect 1406 31445 1432 31509
rect 1496 31445 2700 31509
rect 99 31429 2700 31445
rect 99 31365 982 31429
rect 1046 31365 1072 31429
rect 1136 31365 1162 31429
rect 1226 31365 1252 31429
rect 1316 31365 1342 31429
rect 1406 31365 1432 31429
rect 1496 31365 2700 31429
rect 99 31349 2700 31365
rect 99 31285 982 31349
rect 1046 31285 1072 31349
rect 1136 31285 1162 31349
rect 1226 31285 1252 31349
rect 1316 31285 1342 31349
rect 1406 31285 1432 31349
rect 1496 31285 2700 31349
rect 99 31269 2700 31285
rect 99 31205 982 31269
rect 1046 31205 1072 31269
rect 1136 31205 1162 31269
rect 1226 31205 1252 31269
rect 1316 31205 1342 31269
rect 1406 31205 1432 31269
rect 1496 31205 2700 31269
rect 99 31189 2700 31205
rect 99 31125 982 31189
rect 1046 31125 1072 31189
rect 1136 31125 1162 31189
rect 1226 31125 1252 31189
rect 1316 31125 1342 31189
rect 1406 31125 1432 31189
rect 1496 31125 2700 31189
rect 99 31109 2700 31125
rect 99 31045 982 31109
rect 1046 31045 1072 31109
rect 1136 31045 1162 31109
rect 1226 31045 1252 31109
rect 1316 31045 1342 31109
rect 1406 31045 1432 31109
rect 1496 31045 2700 31109
rect 99 31029 2700 31045
rect 99 30965 982 31029
rect 1046 30965 1072 31029
rect 1136 30965 1162 31029
rect 1226 30965 1252 31029
rect 1316 30965 1342 31029
rect 1406 30965 1432 31029
rect 1496 30965 2700 31029
rect 99 30949 2700 30965
rect 99 30885 982 30949
rect 1046 30885 1072 30949
rect 1136 30885 1162 30949
rect 1226 30885 1252 30949
rect 1316 30885 1342 30949
rect 1406 30885 1432 30949
rect 1496 30885 2700 30949
rect 99 30869 2700 30885
rect 99 30805 982 30869
rect 1046 30805 1072 30869
rect 1136 30805 1162 30869
rect 1226 30805 1252 30869
rect 1316 30805 1342 30869
rect 1406 30805 1432 30869
rect 1496 30805 2700 30869
rect 99 30789 2700 30805
rect 99 30725 982 30789
rect 1046 30725 1072 30789
rect 1136 30725 1162 30789
rect 1226 30725 1252 30789
rect 1316 30725 1342 30789
rect 1406 30725 1432 30789
rect 1496 30725 2700 30789
rect 99 30709 2700 30725
rect 99 30645 982 30709
rect 1046 30645 1072 30709
rect 1136 30645 1162 30709
rect 1226 30645 1252 30709
rect 1316 30645 1342 30709
rect 1406 30645 1432 30709
rect 1496 30645 2700 30709
rect 99 30629 2700 30645
rect 99 30565 982 30629
rect 1046 30565 1072 30629
rect 1136 30565 1162 30629
rect 1226 30565 1252 30629
rect 1316 30565 1342 30629
rect 1406 30565 1432 30629
rect 1496 30565 2700 30629
rect 99 30549 2700 30565
rect 99 30485 982 30549
rect 1046 30485 1072 30549
rect 1136 30485 1162 30549
rect 1226 30485 1252 30549
rect 1316 30485 1342 30549
rect 1406 30485 1432 30549
rect 1496 30485 2700 30549
rect 99 30469 2700 30485
rect 99 30405 982 30469
rect 1046 30405 1072 30469
rect 1136 30405 1162 30469
rect 1226 30405 1252 30469
rect 1316 30405 1342 30469
rect 1406 30405 1432 30469
rect 1496 30405 2700 30469
rect 99 30389 2700 30405
rect 99 30325 982 30389
rect 1046 30325 1072 30389
rect 1136 30325 1162 30389
rect 1226 30325 1252 30389
rect 1316 30325 1342 30389
rect 1406 30325 1432 30389
rect 1496 30325 2700 30389
rect 99 30309 2700 30325
rect 99 30245 982 30309
rect 1046 30245 1072 30309
rect 1136 30245 1162 30309
rect 1226 30245 1252 30309
rect 1316 30245 1342 30309
rect 1406 30245 1432 30309
rect 1496 30245 2700 30309
rect 99 30229 2700 30245
rect 99 30165 982 30229
rect 1046 30165 1072 30229
rect 1136 30165 1162 30229
rect 1226 30165 1252 30229
rect 1316 30165 1342 30229
rect 1406 30165 1432 30229
rect 1496 30165 2700 30229
rect 99 30149 2700 30165
rect 99 30085 982 30149
rect 1046 30085 1072 30149
rect 1136 30085 1162 30149
rect 1226 30085 1252 30149
rect 1316 30085 1342 30149
rect 1406 30085 1432 30149
rect 1496 30085 2700 30149
rect 99 30069 2700 30085
rect 99 30005 982 30069
rect 1046 30005 1072 30069
rect 1136 30005 1162 30069
rect 1226 30005 1252 30069
rect 1316 30005 1342 30069
rect 1406 30005 1432 30069
rect 1496 30005 2700 30069
rect 99 29989 2700 30005
rect 99 29925 982 29989
rect 1046 29925 1072 29989
rect 1136 29925 1162 29989
rect 1226 29925 1252 29989
rect 1316 29925 1342 29989
rect 1406 29925 1432 29989
rect 1496 29925 2700 29989
rect 99 29909 2700 29925
rect 99 29845 982 29909
rect 1046 29845 1072 29909
rect 1136 29845 1162 29909
rect 1226 29845 1252 29909
rect 1316 29845 1342 29909
rect 1406 29845 1432 29909
rect 1496 29845 2700 29909
rect 99 29829 2700 29845
rect 99 29765 982 29829
rect 1046 29765 1072 29829
rect 1136 29765 1162 29829
rect 1226 29765 1252 29829
rect 1316 29765 1342 29829
rect 1406 29765 1432 29829
rect 1496 29765 2700 29829
rect 99 29749 2700 29765
rect 99 29685 982 29749
rect 1046 29685 1072 29749
rect 1136 29685 1162 29749
rect 1226 29685 1252 29749
rect 1316 29685 1342 29749
rect 1406 29685 1432 29749
rect 1496 29685 2700 29749
rect 99 29669 2700 29685
rect 99 29605 982 29669
rect 1046 29605 1072 29669
rect 1136 29605 1162 29669
rect 1226 29605 1252 29669
rect 1316 29605 1342 29669
rect 1406 29605 1432 29669
rect 1496 29605 2700 29669
rect 99 29589 2700 29605
rect 99 29525 982 29589
rect 1046 29525 1072 29589
rect 1136 29525 1162 29589
rect 1226 29525 1252 29589
rect 1316 29525 1342 29589
rect 1406 29525 1432 29589
rect 1496 29525 2700 29589
rect 99 29509 2700 29525
rect 99 29445 982 29509
rect 1046 29445 1072 29509
rect 1136 29445 1162 29509
rect 1226 29445 1252 29509
rect 1316 29445 1342 29509
rect 1406 29445 1432 29509
rect 1496 29445 2700 29509
rect 99 29429 2700 29445
rect 99 29365 982 29429
rect 1046 29365 1072 29429
rect 1136 29365 1162 29429
rect 1226 29365 1252 29429
rect 1316 29365 1342 29429
rect 1406 29365 1432 29429
rect 1496 29365 2700 29429
rect 99 29349 2700 29365
rect 99 29285 982 29349
rect 1046 29285 1072 29349
rect 1136 29285 1162 29349
rect 1226 29285 1252 29349
rect 1316 29285 1342 29349
rect 1406 29285 1432 29349
rect 1496 29285 2700 29349
rect 99 29269 2700 29285
rect 99 29205 982 29269
rect 1046 29205 1072 29269
rect 1136 29205 1162 29269
rect 1226 29205 1252 29269
rect 1316 29205 1342 29269
rect 1406 29205 1432 29269
rect 1496 29205 2700 29269
rect 99 29189 2700 29205
rect 99 29125 982 29189
rect 1046 29125 1072 29189
rect 1136 29125 1162 29189
rect 1226 29125 1252 29189
rect 1316 29125 1342 29189
rect 1406 29125 1432 29189
rect 1496 29125 2700 29189
rect 99 29109 2700 29125
rect 99 29045 982 29109
rect 1046 29045 1072 29109
rect 1136 29045 1162 29109
rect 1226 29045 1252 29109
rect 1316 29045 1342 29109
rect 1406 29045 1432 29109
rect 1496 29045 2700 29109
rect 99 29029 2700 29045
rect 99 28965 982 29029
rect 1046 28965 1072 29029
rect 1136 28965 1162 29029
rect 1226 28965 1252 29029
rect 1316 28965 1342 29029
rect 1406 28965 1432 29029
rect 1496 28965 2700 29029
rect 99 28949 2700 28965
rect 99 28885 982 28949
rect 1046 28885 1072 28949
rect 1136 28885 1162 28949
rect 1226 28885 1252 28949
rect 1316 28885 1342 28949
rect 1406 28885 1432 28949
rect 1496 28885 2700 28949
rect 99 28869 2700 28885
rect 99 28805 982 28869
rect 1046 28805 1072 28869
rect 1136 28805 1162 28869
rect 1226 28805 1252 28869
rect 1316 28805 1342 28869
rect 1406 28805 1432 28869
rect 1496 28805 2700 28869
rect 99 28789 2700 28805
rect 99 28725 982 28789
rect 1046 28725 1072 28789
rect 1136 28725 1162 28789
rect 1226 28725 1252 28789
rect 1316 28725 1342 28789
rect 1406 28725 1432 28789
rect 1496 28725 2700 28789
rect 99 28709 2700 28725
rect 99 28645 982 28709
rect 1046 28645 1072 28709
rect 1136 28645 1162 28709
rect 1226 28645 1252 28709
rect 1316 28645 1342 28709
rect 1406 28645 1432 28709
rect 1496 28645 2700 28709
rect 99 28629 2700 28645
rect 99 28565 982 28629
rect 1046 28565 1072 28629
rect 1136 28565 1162 28629
rect 1226 28565 1252 28629
rect 1316 28565 1342 28629
rect 1406 28565 1432 28629
rect 1496 28565 2700 28629
rect 99 28549 2700 28565
rect 99 28485 982 28549
rect 1046 28485 1072 28549
rect 1136 28485 1162 28549
rect 1226 28485 1252 28549
rect 1316 28485 1342 28549
rect 1406 28485 1432 28549
rect 1496 28485 2700 28549
rect 99 28469 2700 28485
rect 99 28405 982 28469
rect 1046 28405 1072 28469
rect 1136 28405 1162 28469
rect 1226 28405 1252 28469
rect 1316 28405 1342 28469
rect 1406 28405 1432 28469
rect 1496 28405 2700 28469
rect 99 28389 2700 28405
rect 99 28325 982 28389
rect 1046 28325 1072 28389
rect 1136 28325 1162 28389
rect 1226 28325 1252 28389
rect 1316 28325 1342 28389
rect 1406 28325 1432 28389
rect 1496 28325 2700 28389
rect 99 28309 2700 28325
rect 99 28245 982 28309
rect 1046 28245 1072 28309
rect 1136 28245 1162 28309
rect 1226 28245 1252 28309
rect 1316 28245 1342 28309
rect 1406 28245 1432 28309
rect 1496 28245 2700 28309
rect 99 28229 2700 28245
rect 99 28165 982 28229
rect 1046 28165 1072 28229
rect 1136 28165 1162 28229
rect 1226 28165 1252 28229
rect 1316 28165 1342 28229
rect 1406 28165 1432 28229
rect 1496 28165 2700 28229
rect 99 28149 2700 28165
rect 99 28085 982 28149
rect 1046 28085 1072 28149
rect 1136 28085 1162 28149
rect 1226 28085 1252 28149
rect 1316 28085 1342 28149
rect 1406 28085 1432 28149
rect 1496 28085 2700 28149
rect 99 28069 2700 28085
rect 99 28005 982 28069
rect 1046 28005 1072 28069
rect 1136 28005 1162 28069
rect 1226 28005 1252 28069
rect 1316 28005 1342 28069
rect 1406 28005 1432 28069
rect 1496 28005 2700 28069
rect 99 27989 2700 28005
rect 99 27925 982 27989
rect 1046 27925 1072 27989
rect 1136 27925 1162 27989
rect 1226 27925 1252 27989
rect 1316 27925 1342 27989
rect 1406 27925 1432 27989
rect 1496 27925 2700 27989
rect 99 27909 2700 27925
rect 99 27845 982 27909
rect 1046 27845 1072 27909
rect 1136 27845 1162 27909
rect 1226 27845 1252 27909
rect 1316 27845 1342 27909
rect 1406 27845 1432 27909
rect 1496 27845 2700 27909
rect 99 27829 2700 27845
rect 99 27765 982 27829
rect 1046 27765 1072 27829
rect 1136 27765 1162 27829
rect 1226 27765 1252 27829
rect 1316 27765 1342 27829
rect 1406 27765 1432 27829
rect 1496 27765 2700 27829
rect 99 27749 2700 27765
rect 99 27685 982 27749
rect 1046 27685 1072 27749
rect 1136 27685 1162 27749
rect 1226 27685 1252 27749
rect 1316 27685 1342 27749
rect 1406 27685 1432 27749
rect 1496 27685 2700 27749
rect 99 27669 2700 27685
rect 99 27605 982 27669
rect 1046 27605 1072 27669
rect 1136 27605 1162 27669
rect 1226 27605 1252 27669
rect 1316 27605 1342 27669
rect 1406 27605 1432 27669
rect 1496 27605 2700 27669
rect 99 27589 2700 27605
rect 99 27525 982 27589
rect 1046 27525 1072 27589
rect 1136 27525 1162 27589
rect 1226 27525 1252 27589
rect 1316 27525 1342 27589
rect 1406 27525 1432 27589
rect 1496 27525 2700 27589
rect 99 27509 2700 27525
rect 99 27445 982 27509
rect 1046 27445 1072 27509
rect 1136 27445 1162 27509
rect 1226 27445 1252 27509
rect 1316 27445 1342 27509
rect 1406 27445 1432 27509
rect 1496 27445 2700 27509
rect 99 27429 2700 27445
rect 99 27365 982 27429
rect 1046 27365 1072 27429
rect 1136 27365 1162 27429
rect 1226 27365 1252 27429
rect 1316 27365 1342 27429
rect 1406 27365 1432 27429
rect 1496 27365 2700 27429
rect 99 27349 2700 27365
rect 99 27285 982 27349
rect 1046 27285 1072 27349
rect 1136 27285 1162 27349
rect 1226 27285 1252 27349
rect 1316 27285 1342 27349
rect 1406 27285 1432 27349
rect 1496 27285 2700 27349
rect 99 27269 2700 27285
rect 99 27205 982 27269
rect 1046 27205 1072 27269
rect 1136 27205 1162 27269
rect 1226 27205 1252 27269
rect 1316 27205 1342 27269
rect 1406 27205 1432 27269
rect 1496 27205 2700 27269
rect 99 27189 2700 27205
rect 99 27125 982 27189
rect 1046 27125 1072 27189
rect 1136 27125 1162 27189
rect 1226 27125 1252 27189
rect 1316 27125 1342 27189
rect 1406 27125 1432 27189
rect 1496 27125 2700 27189
rect 99 27109 2700 27125
rect 99 27045 982 27109
rect 1046 27045 1072 27109
rect 1136 27045 1162 27109
rect 1226 27045 1252 27109
rect 1316 27045 1342 27109
rect 1406 27045 1432 27109
rect 1496 27045 2700 27109
rect 99 27029 2700 27045
rect 99 26965 982 27029
rect 1046 26965 1072 27029
rect 1136 26965 1162 27029
rect 1226 26965 1252 27029
rect 1316 26965 1342 27029
rect 1406 26965 1432 27029
rect 1496 26965 2700 27029
rect 99 26949 2700 26965
rect 99 26885 982 26949
rect 1046 26885 1072 26949
rect 1136 26885 1162 26949
rect 1226 26885 1252 26949
rect 1316 26885 1342 26949
rect 1406 26885 1432 26949
rect 1496 26885 2700 26949
rect 99 26869 2700 26885
rect 99 26805 982 26869
rect 1046 26805 1072 26869
rect 1136 26805 1162 26869
rect 1226 26805 1252 26869
rect 1316 26805 1342 26869
rect 1406 26805 1432 26869
rect 1496 26805 2700 26869
rect 99 26789 2700 26805
rect 99 26725 982 26789
rect 1046 26725 1072 26789
rect 1136 26725 1162 26789
rect 1226 26725 1252 26789
rect 1316 26725 1342 26789
rect 1406 26725 1432 26789
rect 1496 26725 2700 26789
rect 99 26709 2700 26725
rect 99 26645 982 26709
rect 1046 26645 1072 26709
rect 1136 26645 1162 26709
rect 1226 26645 1252 26709
rect 1316 26645 1342 26709
rect 1406 26645 1432 26709
rect 1496 26645 2700 26709
rect 99 26629 2700 26645
rect 99 26565 982 26629
rect 1046 26565 1072 26629
rect 1136 26565 1162 26629
rect 1226 26565 1252 26629
rect 1316 26565 1342 26629
rect 1406 26565 1432 26629
rect 1496 26565 2700 26629
rect 99 26549 2700 26565
rect 99 26485 982 26549
rect 1046 26485 1072 26549
rect 1136 26485 1162 26549
rect 1226 26485 1252 26549
rect 1316 26485 1342 26549
rect 1406 26485 1432 26549
rect 1496 26485 2700 26549
rect 99 26469 2700 26485
rect 99 26405 982 26469
rect 1046 26405 1072 26469
rect 1136 26405 1162 26469
rect 1226 26405 1252 26469
rect 1316 26405 1342 26469
rect 1406 26405 1432 26469
rect 1496 26405 2700 26469
rect 99 26389 2700 26405
rect 99 26325 982 26389
rect 1046 26325 1072 26389
rect 1136 26325 1162 26389
rect 1226 26325 1252 26389
rect 1316 26325 1342 26389
rect 1406 26325 1432 26389
rect 1496 26325 2700 26389
rect 99 26309 2700 26325
rect 99 26245 982 26309
rect 1046 26245 1072 26309
rect 1136 26245 1162 26309
rect 1226 26245 1252 26309
rect 1316 26245 1342 26309
rect 1406 26245 1432 26309
rect 1496 26245 2700 26309
rect 99 26229 2700 26245
rect 99 26165 982 26229
rect 1046 26165 1072 26229
rect 1136 26165 1162 26229
rect 1226 26165 1252 26229
rect 1316 26165 1342 26229
rect 1406 26165 1432 26229
rect 1496 26165 2700 26229
rect 99 26149 2700 26165
rect 99 26085 982 26149
rect 1046 26085 1072 26149
rect 1136 26085 1162 26149
rect 1226 26085 1252 26149
rect 1316 26085 1342 26149
rect 1406 26085 1432 26149
rect 1496 26085 2700 26149
rect 99 26069 2700 26085
rect 99 26005 982 26069
rect 1046 26005 1072 26069
rect 1136 26005 1162 26069
rect 1226 26005 1252 26069
rect 1316 26005 1342 26069
rect 1406 26005 1432 26069
rect 1496 26005 2700 26069
rect 99 25989 2700 26005
rect 99 25925 982 25989
rect 1046 25925 1072 25989
rect 1136 25925 1162 25989
rect 1226 25925 1252 25989
rect 1316 25925 1342 25989
rect 1406 25925 1432 25989
rect 1496 25925 2700 25989
rect 99 25909 2700 25925
rect 99 25845 982 25909
rect 1046 25845 1072 25909
rect 1136 25845 1162 25909
rect 1226 25845 1252 25909
rect 1316 25845 1342 25909
rect 1406 25845 1432 25909
rect 1496 25845 2700 25909
rect 99 25829 2700 25845
rect 99 25765 982 25829
rect 1046 25765 1072 25829
rect 1136 25765 1162 25829
rect 1226 25765 1252 25829
rect 1316 25765 1342 25829
rect 1406 25765 1432 25829
rect 1496 25765 2700 25829
rect 99 25749 2700 25765
rect 99 25685 982 25749
rect 1046 25685 1072 25749
rect 1136 25685 1162 25749
rect 1226 25685 1252 25749
rect 1316 25685 1342 25749
rect 1406 25685 1432 25749
rect 1496 25685 2700 25749
rect 99 25669 2700 25685
rect 99 25605 982 25669
rect 1046 25605 1072 25669
rect 1136 25605 1162 25669
rect 1226 25605 1252 25669
rect 1316 25605 1342 25669
rect 1406 25605 1432 25669
rect 1496 25605 2700 25669
rect 99 25589 2700 25605
rect 99 25525 982 25589
rect 1046 25525 1072 25589
rect 1136 25525 1162 25589
rect 1226 25525 1252 25589
rect 1316 25525 1342 25589
rect 1406 25525 1432 25589
rect 1496 25525 2700 25589
rect 99 25509 2700 25525
rect 99 25445 982 25509
rect 1046 25445 1072 25509
rect 1136 25445 1162 25509
rect 1226 25445 1252 25509
rect 1316 25445 1342 25509
rect 1406 25445 1432 25509
rect 1496 25445 2700 25509
rect 99 25429 2700 25445
rect 99 25365 982 25429
rect 1046 25365 1072 25429
rect 1136 25365 1162 25429
rect 1226 25365 1252 25429
rect 1316 25365 1342 25429
rect 1406 25365 1432 25429
rect 1496 25365 2700 25429
rect 99 25349 2700 25365
rect 99 25285 982 25349
rect 1046 25285 1072 25349
rect 1136 25285 1162 25349
rect 1226 25285 1252 25349
rect 1316 25285 1342 25349
rect 1406 25285 1432 25349
rect 1496 25285 2700 25349
rect 99 25269 2700 25285
rect 99 25205 982 25269
rect 1046 25205 1072 25269
rect 1136 25205 1162 25269
rect 1226 25205 1252 25269
rect 1316 25205 1342 25269
rect 1406 25205 1432 25269
rect 1496 25205 2700 25269
rect 99 25189 2700 25205
rect 99 25125 982 25189
rect 1046 25125 1072 25189
rect 1136 25125 1162 25189
rect 1226 25125 1252 25189
rect 1316 25125 1342 25189
rect 1406 25125 1432 25189
rect 1496 25125 2700 25189
rect 99 25109 2700 25125
rect 99 25045 982 25109
rect 1046 25045 1072 25109
rect 1136 25045 1162 25109
rect 1226 25045 1252 25109
rect 1316 25045 1342 25109
rect 1406 25045 1432 25109
rect 1496 25045 2700 25109
rect 99 25029 2700 25045
rect 99 24965 982 25029
rect 1046 24965 1072 25029
rect 1136 24965 1162 25029
rect 1226 24965 1252 25029
rect 1316 24965 1342 25029
rect 1406 24965 1432 25029
rect 1496 24965 2700 25029
rect 99 24949 2700 24965
rect 99 24885 982 24949
rect 1046 24885 1072 24949
rect 1136 24885 1162 24949
rect 1226 24885 1252 24949
rect 1316 24885 1342 24949
rect 1406 24885 1432 24949
rect 1496 24885 2700 24949
rect 99 24869 2700 24885
rect 99 24805 982 24869
rect 1046 24805 1072 24869
rect 1136 24805 1162 24869
rect 1226 24805 1252 24869
rect 1316 24805 1342 24869
rect 1406 24805 1432 24869
rect 1496 24805 2700 24869
rect 99 24789 2700 24805
rect 99 24725 982 24789
rect 1046 24725 1072 24789
rect 1136 24725 1162 24789
rect 1226 24725 1252 24789
rect 1316 24725 1342 24789
rect 1406 24725 1432 24789
rect 1496 24725 2700 24789
rect 99 24709 2700 24725
rect 99 24645 982 24709
rect 1046 24645 1072 24709
rect 1136 24645 1162 24709
rect 1226 24645 1252 24709
rect 1316 24645 1342 24709
rect 1406 24645 1432 24709
rect 1496 24645 2700 24709
rect 99 24629 2700 24645
rect 99 24565 982 24629
rect 1046 24565 1072 24629
rect 1136 24565 1162 24629
rect 1226 24565 1252 24629
rect 1316 24565 1342 24629
rect 1406 24565 1432 24629
rect 1496 24565 2700 24629
rect 99 24549 2700 24565
rect 99 24485 982 24549
rect 1046 24485 1072 24549
rect 1136 24485 1162 24549
rect 1226 24485 1252 24549
rect 1316 24485 1342 24549
rect 1406 24485 1432 24549
rect 1496 24485 2700 24549
rect 99 24469 2700 24485
rect 99 24405 982 24469
rect 1046 24405 1072 24469
rect 1136 24405 1162 24469
rect 1226 24405 1252 24469
rect 1316 24405 1342 24469
rect 1406 24405 1432 24469
rect 1496 24405 2700 24469
rect 99 24389 2700 24405
rect 99 24325 982 24389
rect 1046 24325 1072 24389
rect 1136 24325 1162 24389
rect 1226 24325 1252 24389
rect 1316 24325 1342 24389
rect 1406 24325 1432 24389
rect 1496 24325 2700 24389
rect 99 24309 2700 24325
rect 99 24245 982 24309
rect 1046 24245 1072 24309
rect 1136 24245 1162 24309
rect 1226 24245 1252 24309
rect 1316 24245 1342 24309
rect 1406 24245 1432 24309
rect 1496 24245 2700 24309
rect 99 24229 2700 24245
rect 99 24165 982 24229
rect 1046 24165 1072 24229
rect 1136 24165 1162 24229
rect 1226 24165 1252 24229
rect 1316 24165 1342 24229
rect 1406 24165 1432 24229
rect 1496 24165 2700 24229
rect 99 24149 2700 24165
rect 99 24085 982 24149
rect 1046 24085 1072 24149
rect 1136 24085 1162 24149
rect 1226 24085 1252 24149
rect 1316 24085 1342 24149
rect 1406 24085 1432 24149
rect 1496 24085 2700 24149
rect 99 24069 2700 24085
rect 99 24005 982 24069
rect 1046 24005 1072 24069
rect 1136 24005 1162 24069
rect 1226 24005 1252 24069
rect 1316 24005 1342 24069
rect 1406 24005 1432 24069
rect 1496 24005 2700 24069
rect 99 23989 2700 24005
rect 99 23925 982 23989
rect 1046 23925 1072 23989
rect 1136 23925 1162 23989
rect 1226 23925 1252 23989
rect 1316 23925 1342 23989
rect 1406 23925 1432 23989
rect 1496 23925 2700 23989
rect 99 23909 2700 23925
rect 99 23845 982 23909
rect 1046 23845 1072 23909
rect 1136 23845 1162 23909
rect 1226 23845 1252 23909
rect 1316 23845 1342 23909
rect 1406 23845 1432 23909
rect 1496 23845 2700 23909
rect 99 23829 2700 23845
rect 99 23765 982 23829
rect 1046 23765 1072 23829
rect 1136 23765 1162 23829
rect 1226 23765 1252 23829
rect 1316 23765 1342 23829
rect 1406 23765 1432 23829
rect 1496 23765 2700 23829
rect 99 23749 2700 23765
rect 99 23685 982 23749
rect 1046 23685 1072 23749
rect 1136 23685 1162 23749
rect 1226 23685 1252 23749
rect 1316 23685 1342 23749
rect 1406 23685 1432 23749
rect 1496 23685 2700 23749
rect 99 23669 2700 23685
rect 99 23605 982 23669
rect 1046 23605 1072 23669
rect 1136 23605 1162 23669
rect 1226 23605 1252 23669
rect 1316 23605 1342 23669
rect 1406 23605 1432 23669
rect 1496 23605 2700 23669
rect 99 23589 2700 23605
rect 99 23525 982 23589
rect 1046 23525 1072 23589
rect 1136 23525 1162 23589
rect 1226 23525 1252 23589
rect 1316 23525 1342 23589
rect 1406 23525 1432 23589
rect 1496 23525 2700 23589
rect 99 23509 2700 23525
rect 99 23445 982 23509
rect 1046 23445 1072 23509
rect 1136 23445 1162 23509
rect 1226 23445 1252 23509
rect 1316 23445 1342 23509
rect 1406 23445 1432 23509
rect 1496 23445 2700 23509
rect 99 23429 2700 23445
rect 99 23365 982 23429
rect 1046 23365 1072 23429
rect 1136 23365 1162 23429
rect 1226 23365 1252 23429
rect 1316 23365 1342 23429
rect 1406 23365 1432 23429
rect 1496 23365 2700 23429
rect 99 23349 2700 23365
rect 99 23285 982 23349
rect 1046 23285 1072 23349
rect 1136 23285 1162 23349
rect 1226 23285 1252 23349
rect 1316 23285 1342 23349
rect 1406 23285 1432 23349
rect 1496 23285 2700 23349
rect 99 23268 2700 23285
rect 99 23204 982 23268
rect 1046 23204 1072 23268
rect 1136 23204 1162 23268
rect 1226 23204 1252 23268
rect 1316 23204 1342 23268
rect 1406 23204 1432 23268
rect 1496 23204 2700 23268
rect 99 23187 2700 23204
rect 99 23123 982 23187
rect 1046 23123 1072 23187
rect 1136 23123 1162 23187
rect 1226 23123 1252 23187
rect 1316 23123 1342 23187
rect 1406 23123 1432 23187
rect 1496 23123 2700 23187
rect 99 23106 2700 23123
rect 99 23042 982 23106
rect 1046 23042 1072 23106
rect 1136 23042 1162 23106
rect 1226 23042 1252 23106
rect 1316 23042 1342 23106
rect 1406 23042 1432 23106
rect 1496 23042 2700 23106
rect 99 23025 2700 23042
rect 99 22961 982 23025
rect 1046 22961 1072 23025
rect 1136 22961 1162 23025
rect 1226 22961 1252 23025
rect 1316 22961 1342 23025
rect 1406 22961 1432 23025
rect 1496 22961 2700 23025
rect 99 22944 2700 22961
rect 99 22880 982 22944
rect 1046 22880 1072 22944
rect 1136 22880 1162 22944
rect 1226 22880 1252 22944
rect 1316 22880 1342 22944
rect 1406 22880 1432 22944
rect 1496 22880 2700 22944
rect 99 22863 2700 22880
rect 99 22799 982 22863
rect 1046 22799 1072 22863
rect 1136 22799 1162 22863
rect 1226 22799 1252 22863
rect 1316 22799 1342 22863
rect 1406 22799 1432 22863
rect 1496 22799 2700 22863
rect 99 22782 2700 22799
rect 99 22718 982 22782
rect 1046 22718 1072 22782
rect 1136 22718 1162 22782
rect 1226 22718 1252 22782
rect 1316 22718 1342 22782
rect 1406 22718 1432 22782
rect 1496 22718 2700 22782
rect 99 22701 2700 22718
rect 99 22637 982 22701
rect 1046 22637 1072 22701
rect 1136 22637 1162 22701
rect 1226 22637 1252 22701
rect 1316 22637 1342 22701
rect 1406 22637 1432 22701
rect 1496 22637 2700 22701
rect 99 22620 2700 22637
rect 99 22556 982 22620
rect 1046 22556 1072 22620
rect 1136 22556 1162 22620
rect 1226 22556 1252 22620
rect 1316 22556 1342 22620
rect 1406 22556 1432 22620
rect 1496 22556 2700 22620
rect 99 22539 2700 22556
rect 99 22475 982 22539
rect 1046 22475 1072 22539
rect 1136 22475 1162 22539
rect 1226 22475 1252 22539
rect 1316 22475 1342 22539
rect 1406 22475 1432 22539
rect 1496 22475 2700 22539
rect 99 22458 2700 22475
rect 99 22394 982 22458
rect 1046 22394 1072 22458
rect 1136 22394 1162 22458
rect 1226 22394 1252 22458
rect 1316 22394 1342 22458
rect 1406 22394 1432 22458
rect 1496 22394 2700 22458
rect 99 22377 2700 22394
rect 99 22313 982 22377
rect 1046 22313 1072 22377
rect 1136 22313 1162 22377
rect 1226 22313 1252 22377
rect 1316 22313 1342 22377
rect 1406 22313 1432 22377
rect 1496 22313 2700 22377
rect 99 22296 2700 22313
rect 99 22232 982 22296
rect 1046 22232 1072 22296
rect 1136 22232 1162 22296
rect 1226 22232 1252 22296
rect 1316 22232 1342 22296
rect 1406 22232 1432 22296
rect 1496 22232 2700 22296
rect 99 22215 2700 22232
rect 99 22151 982 22215
rect 1046 22151 1072 22215
rect 1136 22151 1162 22215
rect 1226 22151 1252 22215
rect 1316 22151 1342 22215
rect 1406 22151 1432 22215
rect 1496 22151 2700 22215
rect 99 22134 2700 22151
rect 99 22070 982 22134
rect 1046 22070 1072 22134
rect 1136 22070 1162 22134
rect 1226 22070 1252 22134
rect 1316 22070 1342 22134
rect 1406 22070 1432 22134
rect 1496 22070 2700 22134
rect 99 22053 2700 22070
rect 99 21989 982 22053
rect 1046 21989 1072 22053
rect 1136 21989 1162 22053
rect 1226 21989 1252 22053
rect 1316 21989 1342 22053
rect 1406 21989 1432 22053
rect 1496 21989 2700 22053
rect 99 21972 2700 21989
rect 99 21908 982 21972
rect 1046 21908 1072 21972
rect 1136 21908 1162 21972
rect 1226 21908 1252 21972
rect 1316 21908 1342 21972
rect 1406 21908 1432 21972
rect 1496 21908 2700 21972
rect 99 21891 2700 21908
rect 99 21827 982 21891
rect 1046 21827 1072 21891
rect 1136 21827 1162 21891
rect 1226 21827 1252 21891
rect 1316 21827 1342 21891
rect 1406 21827 1432 21891
rect 1496 21827 2700 21891
rect 99 21810 2700 21827
rect 99 21746 982 21810
rect 1046 21746 1072 21810
rect 1136 21746 1162 21810
rect 1226 21746 1252 21810
rect 1316 21746 1342 21810
rect 1406 21746 1432 21810
rect 1496 21746 2700 21810
rect 99 21729 2700 21746
rect 99 21665 982 21729
rect 1046 21665 1072 21729
rect 1136 21665 1162 21729
rect 1226 21665 1252 21729
rect 1316 21665 1342 21729
rect 1406 21665 1432 21729
rect 1496 21665 2700 21729
rect 99 21648 2700 21665
rect 99 21584 982 21648
rect 1046 21584 1072 21648
rect 1136 21584 1162 21648
rect 1226 21584 1252 21648
rect 1316 21584 1342 21648
rect 1406 21584 1432 21648
rect 1496 21584 2700 21648
rect 99 21567 2700 21584
rect 99 21503 982 21567
rect 1046 21503 1072 21567
rect 1136 21503 1162 21567
rect 1226 21503 1252 21567
rect 1316 21503 1342 21567
rect 1406 21503 1432 21567
rect 1496 21503 2700 21567
rect 99 21486 2700 21503
rect 99 21422 982 21486
rect 1046 21422 1072 21486
rect 1136 21422 1162 21486
rect 1226 21422 1252 21486
rect 1316 21422 1342 21486
rect 1406 21422 1432 21486
rect 1496 21422 2700 21486
rect 99 21405 2700 21422
rect 99 21341 982 21405
rect 1046 21341 1072 21405
rect 1136 21341 1162 21405
rect 1226 21341 1252 21405
rect 1316 21341 1342 21405
rect 1406 21341 1432 21405
rect 1496 21341 2700 21405
rect 99 21324 2700 21341
rect 99 21260 982 21324
rect 1046 21260 1072 21324
rect 1136 21260 1162 21324
rect 1226 21260 1252 21324
rect 1316 21260 1342 21324
rect 1406 21260 1432 21324
rect 1496 21260 2700 21324
rect 99 21243 2700 21260
rect 99 21179 982 21243
rect 1046 21179 1072 21243
rect 1136 21179 1162 21243
rect 1226 21179 1252 21243
rect 1316 21179 1342 21243
rect 1406 21179 1432 21243
rect 1496 21179 2700 21243
rect 99 21162 2700 21179
rect 99 21098 982 21162
rect 1046 21098 1072 21162
rect 1136 21098 1162 21162
rect 1226 21098 1252 21162
rect 1316 21098 1342 21162
rect 1406 21098 1432 21162
rect 1496 21098 2700 21162
rect 99 21081 2700 21098
rect 99 21017 982 21081
rect 1046 21017 1072 21081
rect 1136 21017 1162 21081
rect 1226 21017 1252 21081
rect 1316 21017 1342 21081
rect 1406 21017 1432 21081
rect 1496 21017 2700 21081
rect 99 21000 2700 21017
rect 99 20936 982 21000
rect 1046 20936 1072 21000
rect 1136 20936 1162 21000
rect 1226 20936 1252 21000
rect 1316 20936 1342 21000
rect 1406 20936 1432 21000
rect 1496 20939 2700 21000
rect 1496 20936 1531 20939
rect 99 20919 1531 20936
rect 99 20855 982 20919
rect 1046 20855 1072 20919
rect 1136 20855 1162 20919
rect 1226 20855 1252 20919
rect 1316 20855 1342 20919
rect 1406 20855 1432 20919
rect 1496 20875 1531 20919
rect 1595 20875 2700 20939
rect 1496 20855 2700 20875
rect 99 20825 2700 20855
rect 99 20783 1312 20825
rect 99 20719 1141 20783
rect 1205 20761 1312 20783
rect 1376 20761 1401 20825
rect 1465 20761 1491 20825
rect 1555 20761 1581 20825
rect 1645 20761 1671 20825
rect 1735 20761 2700 20825
rect 1205 20719 2700 20761
rect 99 20709 2700 20719
rect 99 20645 1312 20709
rect 1376 20645 1401 20709
rect 1465 20645 1491 20709
rect 1555 20645 1581 20709
rect 1645 20645 1671 20709
rect 1735 20645 2700 20709
rect 99 20631 2700 20645
rect 99 20593 1812 20631
rect 99 20529 1312 20593
rect 1376 20529 1401 20593
rect 1465 20529 1491 20593
rect 1555 20529 1581 20593
rect 1645 20529 1671 20593
rect 1735 20567 1812 20593
rect 1876 20567 2700 20631
rect 1735 20529 2700 20567
rect 99 20505 2700 20529
rect 99 20469 1632 20505
rect 99 20405 1524 20469
rect 1588 20441 1632 20469
rect 1696 20441 1721 20505
rect 1785 20441 1811 20505
rect 1875 20441 1901 20505
rect 1965 20441 1991 20505
rect 2055 20441 2700 20505
rect 1588 20405 2700 20441
rect 99 20389 2700 20405
rect 99 20325 1632 20389
rect 1696 20325 1721 20389
rect 1785 20325 1811 20389
rect 1875 20325 1901 20389
rect 1965 20325 1991 20389
rect 2055 20325 2700 20389
rect 99 20306 2700 20325
rect 99 20273 2137 20306
rect 99 20209 1632 20273
rect 1696 20209 1721 20273
rect 1785 20209 1811 20273
rect 1875 20209 1901 20273
rect 1965 20209 1991 20273
rect 2055 20242 2137 20273
rect 2201 20242 2700 20306
rect 12300 33434 14858 33458
rect 12300 33396 13489 33434
rect 12300 33332 13348 33396
rect 13412 33370 13489 33396
rect 13553 33370 13579 33434
rect 13643 33370 13669 33434
rect 13733 33370 13759 33434
rect 13823 33370 13848 33434
rect 13912 33370 14858 33434
rect 13412 33332 14858 33370
rect 12300 33318 14858 33332
rect 12300 33254 13489 33318
rect 13553 33254 13579 33318
rect 13643 33254 13669 33318
rect 13733 33254 13759 33318
rect 13823 33254 13848 33318
rect 13912 33254 14858 33318
rect 12300 33202 14858 33254
rect 12300 33138 13489 33202
rect 13553 33138 13579 33202
rect 13643 33138 13669 33202
rect 13733 33138 13759 33202
rect 13823 33138 13848 33202
rect 13912 33138 14858 33202
rect 12300 33109 14858 33138
rect 12300 33045 13520 33109
rect 13584 33045 13610 33109
rect 13674 33045 13700 33109
rect 13764 33045 13790 33109
rect 13854 33045 13880 33109
rect 13944 33045 13970 33109
rect 14034 33045 14858 33109
rect 12300 33029 14858 33045
rect 12300 32965 13520 33029
rect 13584 32965 13610 33029
rect 13674 32965 13700 33029
rect 13764 32965 13790 33029
rect 13854 32965 13880 33029
rect 13944 32965 13970 33029
rect 14034 32965 14858 33029
rect 12300 32949 14858 32965
rect 12300 32885 13520 32949
rect 13584 32885 13610 32949
rect 13674 32885 13700 32949
rect 13764 32885 13790 32949
rect 13854 32885 13880 32949
rect 13944 32885 13970 32949
rect 14034 32885 14858 32949
rect 12300 32869 14858 32885
rect 12300 32805 13520 32869
rect 13584 32805 13610 32869
rect 13674 32805 13700 32869
rect 13764 32805 13790 32869
rect 13854 32805 13880 32869
rect 13944 32805 13970 32869
rect 14034 32805 14858 32869
rect 12300 32789 14858 32805
rect 12300 32725 13520 32789
rect 13584 32725 13610 32789
rect 13674 32725 13700 32789
rect 13764 32725 13790 32789
rect 13854 32725 13880 32789
rect 13944 32725 13970 32789
rect 14034 32725 14858 32789
rect 12300 32709 14858 32725
rect 12300 32645 13520 32709
rect 13584 32645 13610 32709
rect 13674 32645 13700 32709
rect 13764 32645 13790 32709
rect 13854 32645 13880 32709
rect 13944 32645 13970 32709
rect 14034 32645 14858 32709
rect 12300 32629 14858 32645
rect 12300 32565 13520 32629
rect 13584 32565 13610 32629
rect 13674 32565 13700 32629
rect 13764 32565 13790 32629
rect 13854 32565 13880 32629
rect 13944 32565 13970 32629
rect 14034 32565 14858 32629
rect 12300 32549 14858 32565
rect 12300 32485 13520 32549
rect 13584 32485 13610 32549
rect 13674 32485 13700 32549
rect 13764 32485 13790 32549
rect 13854 32485 13880 32549
rect 13944 32485 13970 32549
rect 14034 32485 14858 32549
rect 12300 32469 14858 32485
rect 12300 32405 13520 32469
rect 13584 32405 13610 32469
rect 13674 32405 13700 32469
rect 13764 32405 13790 32469
rect 13854 32405 13880 32469
rect 13944 32405 13970 32469
rect 14034 32405 14858 32469
rect 12300 32389 14858 32405
rect 12300 32325 13520 32389
rect 13584 32325 13610 32389
rect 13674 32325 13700 32389
rect 13764 32325 13790 32389
rect 13854 32325 13880 32389
rect 13944 32325 13970 32389
rect 14034 32325 14858 32389
rect 12300 32309 14858 32325
rect 12300 32245 13520 32309
rect 13584 32245 13610 32309
rect 13674 32245 13700 32309
rect 13764 32245 13790 32309
rect 13854 32245 13880 32309
rect 13944 32245 13970 32309
rect 14034 32245 14858 32309
rect 12300 32229 14858 32245
rect 12300 32165 13520 32229
rect 13584 32165 13610 32229
rect 13674 32165 13700 32229
rect 13764 32165 13790 32229
rect 13854 32165 13880 32229
rect 13944 32165 13970 32229
rect 14034 32165 14858 32229
rect 12300 32149 14858 32165
rect 12300 32085 13520 32149
rect 13584 32085 13610 32149
rect 13674 32085 13700 32149
rect 13764 32085 13790 32149
rect 13854 32085 13880 32149
rect 13944 32085 13970 32149
rect 14034 32085 14858 32149
rect 12300 32069 14858 32085
rect 12300 32005 13520 32069
rect 13584 32005 13610 32069
rect 13674 32005 13700 32069
rect 13764 32005 13790 32069
rect 13854 32005 13880 32069
rect 13944 32005 13970 32069
rect 14034 32005 14858 32069
rect 12300 31989 14858 32005
rect 12300 31925 13520 31989
rect 13584 31925 13610 31989
rect 13674 31925 13700 31989
rect 13764 31925 13790 31989
rect 13854 31925 13880 31989
rect 13944 31925 13970 31989
rect 14034 31925 14858 31989
rect 12300 31909 14858 31925
rect 12300 31845 13520 31909
rect 13584 31845 13610 31909
rect 13674 31845 13700 31909
rect 13764 31845 13790 31909
rect 13854 31845 13880 31909
rect 13944 31845 13970 31909
rect 14034 31845 14858 31909
rect 12300 31829 14858 31845
rect 12300 31765 13520 31829
rect 13584 31765 13610 31829
rect 13674 31765 13700 31829
rect 13764 31765 13790 31829
rect 13854 31765 13880 31829
rect 13944 31765 13970 31829
rect 14034 31765 14858 31829
rect 12300 31749 14858 31765
rect 12300 31685 13520 31749
rect 13584 31685 13610 31749
rect 13674 31685 13700 31749
rect 13764 31685 13790 31749
rect 13854 31685 13880 31749
rect 13944 31685 13970 31749
rect 14034 31685 14858 31749
rect 12300 31669 14858 31685
rect 12300 31605 13520 31669
rect 13584 31605 13610 31669
rect 13674 31605 13700 31669
rect 13764 31605 13790 31669
rect 13854 31605 13880 31669
rect 13944 31605 13970 31669
rect 14034 31605 14858 31669
rect 12300 31589 14858 31605
rect 12300 31525 13520 31589
rect 13584 31525 13610 31589
rect 13674 31525 13700 31589
rect 13764 31525 13790 31589
rect 13854 31525 13880 31589
rect 13944 31525 13970 31589
rect 14034 31525 14858 31589
rect 12300 31509 14858 31525
rect 12300 31445 13520 31509
rect 13584 31445 13610 31509
rect 13674 31445 13700 31509
rect 13764 31445 13790 31509
rect 13854 31445 13880 31509
rect 13944 31445 13970 31509
rect 14034 31445 14858 31509
rect 12300 31429 14858 31445
rect 12300 31365 13520 31429
rect 13584 31365 13610 31429
rect 13674 31365 13700 31429
rect 13764 31365 13790 31429
rect 13854 31365 13880 31429
rect 13944 31365 13970 31429
rect 14034 31365 14858 31429
rect 12300 31349 14858 31365
rect 12300 31285 13520 31349
rect 13584 31285 13610 31349
rect 13674 31285 13700 31349
rect 13764 31285 13790 31349
rect 13854 31285 13880 31349
rect 13944 31285 13970 31349
rect 14034 31285 14858 31349
rect 12300 31269 14858 31285
rect 12300 31205 13520 31269
rect 13584 31205 13610 31269
rect 13674 31205 13700 31269
rect 13764 31205 13790 31269
rect 13854 31205 13880 31269
rect 13944 31205 13970 31269
rect 14034 31205 14858 31269
rect 12300 31189 14858 31205
rect 12300 31125 13520 31189
rect 13584 31125 13610 31189
rect 13674 31125 13700 31189
rect 13764 31125 13790 31189
rect 13854 31125 13880 31189
rect 13944 31125 13970 31189
rect 14034 31125 14858 31189
rect 12300 31109 14858 31125
rect 12300 31045 13520 31109
rect 13584 31045 13610 31109
rect 13674 31045 13700 31109
rect 13764 31045 13790 31109
rect 13854 31045 13880 31109
rect 13944 31045 13970 31109
rect 14034 31045 14858 31109
rect 12300 31029 14858 31045
rect 12300 30965 13520 31029
rect 13584 30965 13610 31029
rect 13674 30965 13700 31029
rect 13764 30965 13790 31029
rect 13854 30965 13880 31029
rect 13944 30965 13970 31029
rect 14034 30965 14858 31029
rect 12300 30949 14858 30965
rect 12300 30885 13520 30949
rect 13584 30885 13610 30949
rect 13674 30885 13700 30949
rect 13764 30885 13790 30949
rect 13854 30885 13880 30949
rect 13944 30885 13970 30949
rect 14034 30885 14858 30949
rect 12300 30869 14858 30885
rect 12300 30805 13520 30869
rect 13584 30805 13610 30869
rect 13674 30805 13700 30869
rect 13764 30805 13790 30869
rect 13854 30805 13880 30869
rect 13944 30805 13970 30869
rect 14034 30805 14858 30869
rect 12300 30789 14858 30805
rect 12300 30725 13520 30789
rect 13584 30725 13610 30789
rect 13674 30725 13700 30789
rect 13764 30725 13790 30789
rect 13854 30725 13880 30789
rect 13944 30725 13970 30789
rect 14034 30725 14858 30789
rect 12300 30709 14858 30725
rect 12300 30645 13520 30709
rect 13584 30645 13610 30709
rect 13674 30645 13700 30709
rect 13764 30645 13790 30709
rect 13854 30645 13880 30709
rect 13944 30645 13970 30709
rect 14034 30645 14858 30709
rect 12300 30629 14858 30645
rect 12300 30565 13520 30629
rect 13584 30565 13610 30629
rect 13674 30565 13700 30629
rect 13764 30565 13790 30629
rect 13854 30565 13880 30629
rect 13944 30565 13970 30629
rect 14034 30565 14858 30629
rect 12300 30549 14858 30565
rect 12300 30485 13520 30549
rect 13584 30485 13610 30549
rect 13674 30485 13700 30549
rect 13764 30485 13790 30549
rect 13854 30485 13880 30549
rect 13944 30485 13970 30549
rect 14034 30485 14858 30549
rect 12300 30469 14858 30485
rect 12300 30405 13520 30469
rect 13584 30405 13610 30469
rect 13674 30405 13700 30469
rect 13764 30405 13790 30469
rect 13854 30405 13880 30469
rect 13944 30405 13970 30469
rect 14034 30405 14858 30469
rect 12300 30389 14858 30405
rect 12300 30325 13520 30389
rect 13584 30325 13610 30389
rect 13674 30325 13700 30389
rect 13764 30325 13790 30389
rect 13854 30325 13880 30389
rect 13944 30325 13970 30389
rect 14034 30325 14858 30389
rect 12300 30309 14858 30325
rect 12300 30245 13520 30309
rect 13584 30245 13610 30309
rect 13674 30245 13700 30309
rect 13764 30245 13790 30309
rect 13854 30245 13880 30309
rect 13944 30245 13970 30309
rect 14034 30245 14858 30309
rect 12300 30229 14858 30245
rect 12300 30165 13520 30229
rect 13584 30165 13610 30229
rect 13674 30165 13700 30229
rect 13764 30165 13790 30229
rect 13854 30165 13880 30229
rect 13944 30165 13970 30229
rect 14034 30165 14858 30229
rect 12300 30149 14858 30165
rect 12300 30085 13520 30149
rect 13584 30085 13610 30149
rect 13674 30085 13700 30149
rect 13764 30085 13790 30149
rect 13854 30085 13880 30149
rect 13944 30085 13970 30149
rect 14034 30085 14858 30149
rect 12300 30069 14858 30085
rect 12300 30005 13520 30069
rect 13584 30005 13610 30069
rect 13674 30005 13700 30069
rect 13764 30005 13790 30069
rect 13854 30005 13880 30069
rect 13944 30005 13970 30069
rect 14034 30005 14858 30069
rect 12300 29989 14858 30005
rect 12300 29925 13520 29989
rect 13584 29925 13610 29989
rect 13674 29925 13700 29989
rect 13764 29925 13790 29989
rect 13854 29925 13880 29989
rect 13944 29925 13970 29989
rect 14034 29925 14858 29989
rect 12300 29909 14858 29925
rect 12300 29845 13520 29909
rect 13584 29845 13610 29909
rect 13674 29845 13700 29909
rect 13764 29845 13790 29909
rect 13854 29845 13880 29909
rect 13944 29845 13970 29909
rect 14034 29845 14858 29909
rect 12300 29829 14858 29845
rect 12300 29765 13520 29829
rect 13584 29765 13610 29829
rect 13674 29765 13700 29829
rect 13764 29765 13790 29829
rect 13854 29765 13880 29829
rect 13944 29765 13970 29829
rect 14034 29765 14858 29829
rect 12300 29749 14858 29765
rect 12300 29685 13520 29749
rect 13584 29685 13610 29749
rect 13674 29685 13700 29749
rect 13764 29685 13790 29749
rect 13854 29685 13880 29749
rect 13944 29685 13970 29749
rect 14034 29685 14858 29749
rect 12300 29669 14858 29685
rect 12300 29605 13520 29669
rect 13584 29605 13610 29669
rect 13674 29605 13700 29669
rect 13764 29605 13790 29669
rect 13854 29605 13880 29669
rect 13944 29605 13970 29669
rect 14034 29605 14858 29669
rect 12300 29589 14858 29605
rect 12300 29525 13520 29589
rect 13584 29525 13610 29589
rect 13674 29525 13700 29589
rect 13764 29525 13790 29589
rect 13854 29525 13880 29589
rect 13944 29525 13970 29589
rect 14034 29525 14858 29589
rect 12300 29509 14858 29525
rect 12300 29445 13520 29509
rect 13584 29445 13610 29509
rect 13674 29445 13700 29509
rect 13764 29445 13790 29509
rect 13854 29445 13880 29509
rect 13944 29445 13970 29509
rect 14034 29445 14858 29509
rect 12300 29429 14858 29445
rect 12300 29365 13520 29429
rect 13584 29365 13610 29429
rect 13674 29365 13700 29429
rect 13764 29365 13790 29429
rect 13854 29365 13880 29429
rect 13944 29365 13970 29429
rect 14034 29365 14858 29429
rect 12300 29349 14858 29365
rect 12300 29285 13520 29349
rect 13584 29285 13610 29349
rect 13674 29285 13700 29349
rect 13764 29285 13790 29349
rect 13854 29285 13880 29349
rect 13944 29285 13970 29349
rect 14034 29285 14858 29349
rect 12300 29269 14858 29285
rect 12300 29205 13520 29269
rect 13584 29205 13610 29269
rect 13674 29205 13700 29269
rect 13764 29205 13790 29269
rect 13854 29205 13880 29269
rect 13944 29205 13970 29269
rect 14034 29205 14858 29269
rect 12300 29189 14858 29205
rect 12300 29125 13520 29189
rect 13584 29125 13610 29189
rect 13674 29125 13700 29189
rect 13764 29125 13790 29189
rect 13854 29125 13880 29189
rect 13944 29125 13970 29189
rect 14034 29125 14858 29189
rect 12300 29109 14858 29125
rect 12300 29045 13520 29109
rect 13584 29045 13610 29109
rect 13674 29045 13700 29109
rect 13764 29045 13790 29109
rect 13854 29045 13880 29109
rect 13944 29045 13970 29109
rect 14034 29045 14858 29109
rect 12300 29029 14858 29045
rect 12300 28965 13520 29029
rect 13584 28965 13610 29029
rect 13674 28965 13700 29029
rect 13764 28965 13790 29029
rect 13854 28965 13880 29029
rect 13944 28965 13970 29029
rect 14034 28965 14858 29029
rect 12300 28949 14858 28965
rect 12300 28885 13520 28949
rect 13584 28885 13610 28949
rect 13674 28885 13700 28949
rect 13764 28885 13790 28949
rect 13854 28885 13880 28949
rect 13944 28885 13970 28949
rect 14034 28885 14858 28949
rect 12300 28869 14858 28885
rect 12300 28805 13520 28869
rect 13584 28805 13610 28869
rect 13674 28805 13700 28869
rect 13764 28805 13790 28869
rect 13854 28805 13880 28869
rect 13944 28805 13970 28869
rect 14034 28805 14858 28869
rect 12300 28789 14858 28805
rect 12300 28725 13520 28789
rect 13584 28725 13610 28789
rect 13674 28725 13700 28789
rect 13764 28725 13790 28789
rect 13854 28725 13880 28789
rect 13944 28725 13970 28789
rect 14034 28725 14858 28789
rect 12300 28709 14858 28725
rect 12300 28645 13520 28709
rect 13584 28645 13610 28709
rect 13674 28645 13700 28709
rect 13764 28645 13790 28709
rect 13854 28645 13880 28709
rect 13944 28645 13970 28709
rect 14034 28645 14858 28709
rect 12300 28629 14858 28645
rect 12300 28565 13520 28629
rect 13584 28565 13610 28629
rect 13674 28565 13700 28629
rect 13764 28565 13790 28629
rect 13854 28565 13880 28629
rect 13944 28565 13970 28629
rect 14034 28565 14858 28629
rect 12300 28549 14858 28565
rect 12300 28485 13520 28549
rect 13584 28485 13610 28549
rect 13674 28485 13700 28549
rect 13764 28485 13790 28549
rect 13854 28485 13880 28549
rect 13944 28485 13970 28549
rect 14034 28485 14858 28549
rect 12300 28469 14858 28485
rect 12300 28405 13520 28469
rect 13584 28405 13610 28469
rect 13674 28405 13700 28469
rect 13764 28405 13790 28469
rect 13854 28405 13880 28469
rect 13944 28405 13970 28469
rect 14034 28405 14858 28469
rect 12300 28389 14858 28405
rect 12300 28325 13520 28389
rect 13584 28325 13610 28389
rect 13674 28325 13700 28389
rect 13764 28325 13790 28389
rect 13854 28325 13880 28389
rect 13944 28325 13970 28389
rect 14034 28325 14858 28389
rect 12300 28309 14858 28325
rect 12300 28245 13520 28309
rect 13584 28245 13610 28309
rect 13674 28245 13700 28309
rect 13764 28245 13790 28309
rect 13854 28245 13880 28309
rect 13944 28245 13970 28309
rect 14034 28245 14858 28309
rect 12300 28229 14858 28245
rect 12300 28165 13520 28229
rect 13584 28165 13610 28229
rect 13674 28165 13700 28229
rect 13764 28165 13790 28229
rect 13854 28165 13880 28229
rect 13944 28165 13970 28229
rect 14034 28165 14858 28229
rect 12300 28149 14858 28165
rect 12300 28085 13520 28149
rect 13584 28085 13610 28149
rect 13674 28085 13700 28149
rect 13764 28085 13790 28149
rect 13854 28085 13880 28149
rect 13944 28085 13970 28149
rect 14034 28085 14858 28149
rect 12300 28069 14858 28085
rect 12300 28005 13520 28069
rect 13584 28005 13610 28069
rect 13674 28005 13700 28069
rect 13764 28005 13790 28069
rect 13854 28005 13880 28069
rect 13944 28005 13970 28069
rect 14034 28005 14858 28069
rect 12300 27989 14858 28005
rect 12300 27925 13520 27989
rect 13584 27925 13610 27989
rect 13674 27925 13700 27989
rect 13764 27925 13790 27989
rect 13854 27925 13880 27989
rect 13944 27925 13970 27989
rect 14034 27925 14858 27989
rect 12300 27909 14858 27925
rect 12300 27845 13520 27909
rect 13584 27845 13610 27909
rect 13674 27845 13700 27909
rect 13764 27845 13790 27909
rect 13854 27845 13880 27909
rect 13944 27845 13970 27909
rect 14034 27845 14858 27909
rect 12300 27829 14858 27845
rect 12300 27765 13520 27829
rect 13584 27765 13610 27829
rect 13674 27765 13700 27829
rect 13764 27765 13790 27829
rect 13854 27765 13880 27829
rect 13944 27765 13970 27829
rect 14034 27765 14858 27829
rect 12300 27749 14858 27765
rect 12300 27685 13520 27749
rect 13584 27685 13610 27749
rect 13674 27685 13700 27749
rect 13764 27685 13790 27749
rect 13854 27685 13880 27749
rect 13944 27685 13970 27749
rect 14034 27685 14858 27749
rect 12300 27669 14858 27685
rect 12300 27605 13520 27669
rect 13584 27605 13610 27669
rect 13674 27605 13700 27669
rect 13764 27605 13790 27669
rect 13854 27605 13880 27669
rect 13944 27605 13970 27669
rect 14034 27605 14858 27669
rect 12300 27589 14858 27605
rect 12300 27525 13520 27589
rect 13584 27525 13610 27589
rect 13674 27525 13700 27589
rect 13764 27525 13790 27589
rect 13854 27525 13880 27589
rect 13944 27525 13970 27589
rect 14034 27525 14858 27589
rect 12300 27509 14858 27525
rect 12300 27445 13520 27509
rect 13584 27445 13610 27509
rect 13674 27445 13700 27509
rect 13764 27445 13790 27509
rect 13854 27445 13880 27509
rect 13944 27445 13970 27509
rect 14034 27445 14858 27509
rect 12300 27429 14858 27445
rect 12300 27365 13520 27429
rect 13584 27365 13610 27429
rect 13674 27365 13700 27429
rect 13764 27365 13790 27429
rect 13854 27365 13880 27429
rect 13944 27365 13970 27429
rect 14034 27365 14858 27429
rect 12300 27349 14858 27365
rect 12300 27285 13520 27349
rect 13584 27285 13610 27349
rect 13674 27285 13700 27349
rect 13764 27285 13790 27349
rect 13854 27285 13880 27349
rect 13944 27285 13970 27349
rect 14034 27285 14858 27349
rect 12300 27269 14858 27285
rect 12300 27205 13520 27269
rect 13584 27205 13610 27269
rect 13674 27205 13700 27269
rect 13764 27205 13790 27269
rect 13854 27205 13880 27269
rect 13944 27205 13970 27269
rect 14034 27205 14858 27269
rect 12300 27189 14858 27205
rect 12300 27125 13520 27189
rect 13584 27125 13610 27189
rect 13674 27125 13700 27189
rect 13764 27125 13790 27189
rect 13854 27125 13880 27189
rect 13944 27125 13970 27189
rect 14034 27125 14858 27189
rect 12300 27109 14858 27125
rect 12300 27045 13520 27109
rect 13584 27045 13610 27109
rect 13674 27045 13700 27109
rect 13764 27045 13790 27109
rect 13854 27045 13880 27109
rect 13944 27045 13970 27109
rect 14034 27045 14858 27109
rect 12300 27029 14858 27045
rect 12300 26965 13520 27029
rect 13584 26965 13610 27029
rect 13674 26965 13700 27029
rect 13764 26965 13790 27029
rect 13854 26965 13880 27029
rect 13944 26965 13970 27029
rect 14034 26965 14858 27029
rect 12300 26949 14858 26965
rect 12300 26885 13520 26949
rect 13584 26885 13610 26949
rect 13674 26885 13700 26949
rect 13764 26885 13790 26949
rect 13854 26885 13880 26949
rect 13944 26885 13970 26949
rect 14034 26885 14858 26949
rect 12300 26869 14858 26885
rect 12300 26805 13520 26869
rect 13584 26805 13610 26869
rect 13674 26805 13700 26869
rect 13764 26805 13790 26869
rect 13854 26805 13880 26869
rect 13944 26805 13970 26869
rect 14034 26805 14858 26869
rect 12300 26789 14858 26805
rect 12300 26725 13520 26789
rect 13584 26725 13610 26789
rect 13674 26725 13700 26789
rect 13764 26725 13790 26789
rect 13854 26725 13880 26789
rect 13944 26725 13970 26789
rect 14034 26725 14858 26789
rect 12300 26709 14858 26725
rect 12300 26645 13520 26709
rect 13584 26645 13610 26709
rect 13674 26645 13700 26709
rect 13764 26645 13790 26709
rect 13854 26645 13880 26709
rect 13944 26645 13970 26709
rect 14034 26645 14858 26709
rect 12300 26629 14858 26645
rect 12300 26565 13520 26629
rect 13584 26565 13610 26629
rect 13674 26565 13700 26629
rect 13764 26565 13790 26629
rect 13854 26565 13880 26629
rect 13944 26565 13970 26629
rect 14034 26565 14858 26629
rect 12300 26549 14858 26565
rect 12300 26485 13520 26549
rect 13584 26485 13610 26549
rect 13674 26485 13700 26549
rect 13764 26485 13790 26549
rect 13854 26485 13880 26549
rect 13944 26485 13970 26549
rect 14034 26485 14858 26549
rect 12300 26469 14858 26485
rect 12300 26405 13520 26469
rect 13584 26405 13610 26469
rect 13674 26405 13700 26469
rect 13764 26405 13790 26469
rect 13854 26405 13880 26469
rect 13944 26405 13970 26469
rect 14034 26405 14858 26469
rect 12300 26389 14858 26405
rect 12300 26325 13520 26389
rect 13584 26325 13610 26389
rect 13674 26325 13700 26389
rect 13764 26325 13790 26389
rect 13854 26325 13880 26389
rect 13944 26325 13970 26389
rect 14034 26325 14858 26389
rect 12300 26309 14858 26325
rect 12300 26245 13520 26309
rect 13584 26245 13610 26309
rect 13674 26245 13700 26309
rect 13764 26245 13790 26309
rect 13854 26245 13880 26309
rect 13944 26245 13970 26309
rect 14034 26245 14858 26309
rect 12300 26229 14858 26245
rect 12300 26165 13520 26229
rect 13584 26165 13610 26229
rect 13674 26165 13700 26229
rect 13764 26165 13790 26229
rect 13854 26165 13880 26229
rect 13944 26165 13970 26229
rect 14034 26165 14858 26229
rect 12300 26149 14858 26165
rect 12300 26085 13520 26149
rect 13584 26085 13610 26149
rect 13674 26085 13700 26149
rect 13764 26085 13790 26149
rect 13854 26085 13880 26149
rect 13944 26085 13970 26149
rect 14034 26085 14858 26149
rect 12300 26069 14858 26085
rect 12300 26005 13520 26069
rect 13584 26005 13610 26069
rect 13674 26005 13700 26069
rect 13764 26005 13790 26069
rect 13854 26005 13880 26069
rect 13944 26005 13970 26069
rect 14034 26005 14858 26069
rect 12300 25989 14858 26005
rect 12300 25925 13520 25989
rect 13584 25925 13610 25989
rect 13674 25925 13700 25989
rect 13764 25925 13790 25989
rect 13854 25925 13880 25989
rect 13944 25925 13970 25989
rect 14034 25925 14858 25989
rect 12300 25909 14858 25925
rect 12300 25845 13520 25909
rect 13584 25845 13610 25909
rect 13674 25845 13700 25909
rect 13764 25845 13790 25909
rect 13854 25845 13880 25909
rect 13944 25845 13970 25909
rect 14034 25845 14858 25909
rect 12300 25829 14858 25845
rect 12300 25765 13520 25829
rect 13584 25765 13610 25829
rect 13674 25765 13700 25829
rect 13764 25765 13790 25829
rect 13854 25765 13880 25829
rect 13944 25765 13970 25829
rect 14034 25765 14858 25829
rect 12300 25749 14858 25765
rect 12300 25685 13520 25749
rect 13584 25685 13610 25749
rect 13674 25685 13700 25749
rect 13764 25685 13790 25749
rect 13854 25685 13880 25749
rect 13944 25685 13970 25749
rect 14034 25685 14858 25749
rect 12300 25669 14858 25685
rect 12300 25605 13520 25669
rect 13584 25605 13610 25669
rect 13674 25605 13700 25669
rect 13764 25605 13790 25669
rect 13854 25605 13880 25669
rect 13944 25605 13970 25669
rect 14034 25605 14858 25669
rect 12300 25589 14858 25605
rect 12300 25525 13520 25589
rect 13584 25525 13610 25589
rect 13674 25525 13700 25589
rect 13764 25525 13790 25589
rect 13854 25525 13880 25589
rect 13944 25525 13970 25589
rect 14034 25525 14858 25589
rect 12300 25509 14858 25525
rect 12300 25445 13520 25509
rect 13584 25445 13610 25509
rect 13674 25445 13700 25509
rect 13764 25445 13790 25509
rect 13854 25445 13880 25509
rect 13944 25445 13970 25509
rect 14034 25445 14858 25509
rect 12300 25429 14858 25445
rect 12300 25365 13520 25429
rect 13584 25365 13610 25429
rect 13674 25365 13700 25429
rect 13764 25365 13790 25429
rect 13854 25365 13880 25429
rect 13944 25365 13970 25429
rect 14034 25365 14858 25429
rect 12300 25349 14858 25365
rect 12300 25285 13520 25349
rect 13584 25285 13610 25349
rect 13674 25285 13700 25349
rect 13764 25285 13790 25349
rect 13854 25285 13880 25349
rect 13944 25285 13970 25349
rect 14034 25285 14858 25349
rect 12300 25269 14858 25285
rect 12300 25205 13520 25269
rect 13584 25205 13610 25269
rect 13674 25205 13700 25269
rect 13764 25205 13790 25269
rect 13854 25205 13880 25269
rect 13944 25205 13970 25269
rect 14034 25205 14858 25269
rect 12300 25189 14858 25205
rect 12300 25125 13520 25189
rect 13584 25125 13610 25189
rect 13674 25125 13700 25189
rect 13764 25125 13790 25189
rect 13854 25125 13880 25189
rect 13944 25125 13970 25189
rect 14034 25125 14858 25189
rect 12300 25109 14858 25125
rect 12300 25045 13520 25109
rect 13584 25045 13610 25109
rect 13674 25045 13700 25109
rect 13764 25045 13790 25109
rect 13854 25045 13880 25109
rect 13944 25045 13970 25109
rect 14034 25045 14858 25109
rect 12300 25029 14858 25045
rect 12300 24965 13520 25029
rect 13584 24965 13610 25029
rect 13674 24965 13700 25029
rect 13764 24965 13790 25029
rect 13854 24965 13880 25029
rect 13944 24965 13970 25029
rect 14034 24965 14858 25029
rect 12300 24949 14858 24965
rect 12300 24885 13520 24949
rect 13584 24885 13610 24949
rect 13674 24885 13700 24949
rect 13764 24885 13790 24949
rect 13854 24885 13880 24949
rect 13944 24885 13970 24949
rect 14034 24885 14858 24949
rect 12300 24869 14858 24885
rect 12300 24805 13520 24869
rect 13584 24805 13610 24869
rect 13674 24805 13700 24869
rect 13764 24805 13790 24869
rect 13854 24805 13880 24869
rect 13944 24805 13970 24869
rect 14034 24805 14858 24869
rect 12300 24789 14858 24805
rect 12300 24725 13520 24789
rect 13584 24725 13610 24789
rect 13674 24725 13700 24789
rect 13764 24725 13790 24789
rect 13854 24725 13880 24789
rect 13944 24725 13970 24789
rect 14034 24725 14858 24789
rect 12300 24709 14858 24725
rect 12300 24645 13520 24709
rect 13584 24645 13610 24709
rect 13674 24645 13700 24709
rect 13764 24645 13790 24709
rect 13854 24645 13880 24709
rect 13944 24645 13970 24709
rect 14034 24645 14858 24709
rect 12300 24629 14858 24645
rect 12300 24565 13520 24629
rect 13584 24565 13610 24629
rect 13674 24565 13700 24629
rect 13764 24565 13790 24629
rect 13854 24565 13880 24629
rect 13944 24565 13970 24629
rect 14034 24565 14858 24629
rect 12300 24549 14858 24565
rect 12300 24485 13520 24549
rect 13584 24485 13610 24549
rect 13674 24485 13700 24549
rect 13764 24485 13790 24549
rect 13854 24485 13880 24549
rect 13944 24485 13970 24549
rect 14034 24485 14858 24549
rect 12300 24469 14858 24485
rect 12300 24405 13520 24469
rect 13584 24405 13610 24469
rect 13674 24405 13700 24469
rect 13764 24405 13790 24469
rect 13854 24405 13880 24469
rect 13944 24405 13970 24469
rect 14034 24405 14858 24469
rect 12300 24389 14858 24405
rect 12300 24325 13520 24389
rect 13584 24325 13610 24389
rect 13674 24325 13700 24389
rect 13764 24325 13790 24389
rect 13854 24325 13880 24389
rect 13944 24325 13970 24389
rect 14034 24325 14858 24389
rect 12300 24309 14858 24325
rect 12300 24245 13520 24309
rect 13584 24245 13610 24309
rect 13674 24245 13700 24309
rect 13764 24245 13790 24309
rect 13854 24245 13880 24309
rect 13944 24245 13970 24309
rect 14034 24245 14858 24309
rect 12300 24229 14858 24245
rect 12300 24165 13520 24229
rect 13584 24165 13610 24229
rect 13674 24165 13700 24229
rect 13764 24165 13790 24229
rect 13854 24165 13880 24229
rect 13944 24165 13970 24229
rect 14034 24165 14858 24229
rect 12300 24149 14858 24165
rect 12300 24085 13520 24149
rect 13584 24085 13610 24149
rect 13674 24085 13700 24149
rect 13764 24085 13790 24149
rect 13854 24085 13880 24149
rect 13944 24085 13970 24149
rect 14034 24085 14858 24149
rect 12300 24069 14858 24085
rect 12300 24005 13520 24069
rect 13584 24005 13610 24069
rect 13674 24005 13700 24069
rect 13764 24005 13790 24069
rect 13854 24005 13880 24069
rect 13944 24005 13970 24069
rect 14034 24005 14858 24069
rect 12300 23989 14858 24005
rect 12300 23925 13520 23989
rect 13584 23925 13610 23989
rect 13674 23925 13700 23989
rect 13764 23925 13790 23989
rect 13854 23925 13880 23989
rect 13944 23925 13970 23989
rect 14034 23925 14858 23989
rect 12300 23909 14858 23925
rect 12300 23845 13520 23909
rect 13584 23845 13610 23909
rect 13674 23845 13700 23909
rect 13764 23845 13790 23909
rect 13854 23845 13880 23909
rect 13944 23845 13970 23909
rect 14034 23845 14858 23909
rect 12300 23829 14858 23845
rect 12300 23765 13520 23829
rect 13584 23765 13610 23829
rect 13674 23765 13700 23829
rect 13764 23765 13790 23829
rect 13854 23765 13880 23829
rect 13944 23765 13970 23829
rect 14034 23765 14858 23829
rect 12300 23749 14858 23765
rect 12300 23685 13520 23749
rect 13584 23685 13610 23749
rect 13674 23685 13700 23749
rect 13764 23685 13790 23749
rect 13854 23685 13880 23749
rect 13944 23685 13970 23749
rect 14034 23685 14858 23749
rect 12300 23669 14858 23685
rect 12300 23605 13520 23669
rect 13584 23605 13610 23669
rect 13674 23605 13700 23669
rect 13764 23605 13790 23669
rect 13854 23605 13880 23669
rect 13944 23605 13970 23669
rect 14034 23605 14858 23669
rect 12300 23589 14858 23605
rect 12300 23525 13520 23589
rect 13584 23525 13610 23589
rect 13674 23525 13700 23589
rect 13764 23525 13790 23589
rect 13854 23525 13880 23589
rect 13944 23525 13970 23589
rect 14034 23525 14858 23589
rect 12300 23509 14858 23525
rect 12300 23445 13520 23509
rect 13584 23445 13610 23509
rect 13674 23445 13700 23509
rect 13764 23445 13790 23509
rect 13854 23445 13880 23509
rect 13944 23445 13970 23509
rect 14034 23445 14858 23509
rect 12300 23429 14858 23445
rect 12300 23365 13520 23429
rect 13584 23365 13610 23429
rect 13674 23365 13700 23429
rect 13764 23365 13790 23429
rect 13854 23365 13880 23429
rect 13944 23365 13970 23429
rect 14034 23365 14858 23429
rect 12300 23349 14858 23365
rect 12300 23285 13520 23349
rect 13584 23285 13610 23349
rect 13674 23285 13700 23349
rect 13764 23285 13790 23349
rect 13854 23285 13880 23349
rect 13944 23285 13970 23349
rect 14034 23285 14858 23349
rect 12300 23268 14858 23285
rect 12300 23204 13520 23268
rect 13584 23204 13610 23268
rect 13674 23204 13700 23268
rect 13764 23204 13790 23268
rect 13854 23204 13880 23268
rect 13944 23204 13970 23268
rect 14034 23204 14858 23268
rect 12300 23187 14858 23204
rect 12300 23123 13520 23187
rect 13584 23123 13610 23187
rect 13674 23123 13700 23187
rect 13764 23123 13790 23187
rect 13854 23123 13880 23187
rect 13944 23123 13970 23187
rect 14034 23123 14858 23187
rect 12300 23106 14858 23123
rect 12300 23042 13520 23106
rect 13584 23042 13610 23106
rect 13674 23042 13700 23106
rect 13764 23042 13790 23106
rect 13854 23042 13880 23106
rect 13944 23042 13970 23106
rect 14034 23042 14858 23106
rect 12300 23025 14858 23042
rect 12300 22961 13520 23025
rect 13584 22961 13610 23025
rect 13674 22961 13700 23025
rect 13764 22961 13790 23025
rect 13854 22961 13880 23025
rect 13944 22961 13970 23025
rect 14034 22961 14858 23025
rect 12300 22944 14858 22961
rect 12300 22880 13520 22944
rect 13584 22880 13610 22944
rect 13674 22880 13700 22944
rect 13764 22880 13790 22944
rect 13854 22880 13880 22944
rect 13944 22880 13970 22944
rect 14034 22880 14858 22944
rect 12300 22863 14858 22880
rect 12300 22799 13520 22863
rect 13584 22799 13610 22863
rect 13674 22799 13700 22863
rect 13764 22799 13790 22863
rect 13854 22799 13880 22863
rect 13944 22799 13970 22863
rect 14034 22799 14858 22863
rect 12300 22782 14858 22799
rect 12300 22718 13520 22782
rect 13584 22718 13610 22782
rect 13674 22718 13700 22782
rect 13764 22718 13790 22782
rect 13854 22718 13880 22782
rect 13944 22718 13970 22782
rect 14034 22718 14858 22782
rect 12300 22701 14858 22718
rect 12300 22637 13520 22701
rect 13584 22637 13610 22701
rect 13674 22637 13700 22701
rect 13764 22637 13790 22701
rect 13854 22637 13880 22701
rect 13944 22637 13970 22701
rect 14034 22637 14858 22701
rect 12300 22620 14858 22637
rect 12300 22556 13520 22620
rect 13584 22556 13610 22620
rect 13674 22556 13700 22620
rect 13764 22556 13790 22620
rect 13854 22556 13880 22620
rect 13944 22556 13970 22620
rect 14034 22556 14858 22620
rect 12300 22539 14858 22556
rect 12300 22475 13520 22539
rect 13584 22475 13610 22539
rect 13674 22475 13700 22539
rect 13764 22475 13790 22539
rect 13854 22475 13880 22539
rect 13944 22475 13970 22539
rect 14034 22475 14858 22539
rect 12300 22458 14858 22475
rect 12300 22394 13520 22458
rect 13584 22394 13610 22458
rect 13674 22394 13700 22458
rect 13764 22394 13790 22458
rect 13854 22394 13880 22458
rect 13944 22394 13970 22458
rect 14034 22394 14858 22458
rect 12300 22377 14858 22394
rect 12300 22313 13520 22377
rect 13584 22313 13610 22377
rect 13674 22313 13700 22377
rect 13764 22313 13790 22377
rect 13854 22313 13880 22377
rect 13944 22313 13970 22377
rect 14034 22313 14858 22377
rect 12300 22296 14858 22313
rect 12300 22232 13520 22296
rect 13584 22232 13610 22296
rect 13674 22232 13700 22296
rect 13764 22232 13790 22296
rect 13854 22232 13880 22296
rect 13944 22232 13970 22296
rect 14034 22232 14858 22296
rect 12300 22215 14858 22232
rect 12300 22151 13520 22215
rect 13584 22151 13610 22215
rect 13674 22151 13700 22215
rect 13764 22151 13790 22215
rect 13854 22151 13880 22215
rect 13944 22151 13970 22215
rect 14034 22151 14858 22215
rect 12300 22134 14858 22151
rect 12300 22070 13520 22134
rect 13584 22070 13610 22134
rect 13674 22070 13700 22134
rect 13764 22070 13790 22134
rect 13854 22070 13880 22134
rect 13944 22070 13970 22134
rect 14034 22070 14858 22134
rect 12300 22053 14858 22070
rect 12300 21989 13520 22053
rect 13584 21989 13610 22053
rect 13674 21989 13700 22053
rect 13764 21989 13790 22053
rect 13854 21989 13880 22053
rect 13944 21989 13970 22053
rect 14034 21989 14858 22053
rect 12300 21972 14858 21989
rect 12300 21908 13520 21972
rect 13584 21908 13610 21972
rect 13674 21908 13700 21972
rect 13764 21908 13790 21972
rect 13854 21908 13880 21972
rect 13944 21908 13970 21972
rect 14034 21908 14858 21972
rect 12300 21891 14858 21908
rect 12300 21827 13520 21891
rect 13584 21827 13610 21891
rect 13674 21827 13700 21891
rect 13764 21827 13790 21891
rect 13854 21827 13880 21891
rect 13944 21827 13970 21891
rect 14034 21827 14858 21891
rect 12300 21810 14858 21827
rect 12300 21746 13520 21810
rect 13584 21746 13610 21810
rect 13674 21746 13700 21810
rect 13764 21746 13790 21810
rect 13854 21746 13880 21810
rect 13944 21746 13970 21810
rect 14034 21746 14858 21810
rect 12300 21729 14858 21746
rect 12300 21665 13520 21729
rect 13584 21665 13610 21729
rect 13674 21665 13700 21729
rect 13764 21665 13790 21729
rect 13854 21665 13880 21729
rect 13944 21665 13970 21729
rect 14034 21665 14858 21729
rect 12300 21648 14858 21665
rect 12300 21584 13520 21648
rect 13584 21584 13610 21648
rect 13674 21584 13700 21648
rect 13764 21584 13790 21648
rect 13854 21584 13880 21648
rect 13944 21584 13970 21648
rect 14034 21584 14858 21648
rect 12300 21567 14858 21584
rect 12300 21503 13520 21567
rect 13584 21503 13610 21567
rect 13674 21503 13700 21567
rect 13764 21503 13790 21567
rect 13854 21503 13880 21567
rect 13944 21503 13970 21567
rect 14034 21503 14858 21567
rect 12300 21486 14858 21503
rect 12300 21422 13520 21486
rect 13584 21422 13610 21486
rect 13674 21422 13700 21486
rect 13764 21422 13790 21486
rect 13854 21422 13880 21486
rect 13944 21422 13970 21486
rect 14034 21422 14858 21486
rect 12300 21405 14858 21422
rect 12300 21341 13520 21405
rect 13584 21341 13610 21405
rect 13674 21341 13700 21405
rect 13764 21341 13790 21405
rect 13854 21341 13880 21405
rect 13944 21341 13970 21405
rect 14034 21341 14858 21405
rect 12300 21324 14858 21341
rect 12300 21260 13520 21324
rect 13584 21260 13610 21324
rect 13674 21260 13700 21324
rect 13764 21260 13790 21324
rect 13854 21260 13880 21324
rect 13944 21260 13970 21324
rect 14034 21260 14858 21324
rect 12300 21243 14858 21260
rect 12300 21179 13520 21243
rect 13584 21179 13610 21243
rect 13674 21179 13700 21243
rect 13764 21179 13790 21243
rect 13854 21179 13880 21243
rect 13944 21179 13970 21243
rect 14034 21179 14858 21243
rect 12300 21162 14858 21179
rect 12300 21098 13520 21162
rect 13584 21098 13610 21162
rect 13674 21098 13700 21162
rect 13764 21098 13790 21162
rect 13854 21098 13880 21162
rect 13944 21098 13970 21162
rect 14034 21098 14858 21162
rect 12300 21081 14858 21098
rect 12300 21017 13520 21081
rect 13584 21017 13610 21081
rect 13674 21017 13700 21081
rect 13764 21017 13790 21081
rect 13854 21017 13880 21081
rect 13944 21017 13970 21081
rect 14034 21017 14858 21081
rect 12300 21000 14858 21017
rect 12300 20939 13520 21000
rect 12300 20875 13421 20939
rect 13485 20936 13520 20939
rect 13584 20936 13610 21000
rect 13674 20936 13700 21000
rect 13764 20936 13790 21000
rect 13854 20936 13880 21000
rect 13944 20936 13970 21000
rect 14034 20936 14858 21000
rect 13485 20919 14858 20936
rect 13485 20875 13520 20919
rect 12300 20855 13520 20875
rect 13584 20855 13610 20919
rect 13674 20855 13700 20919
rect 13764 20855 13790 20919
rect 13854 20855 13880 20919
rect 13944 20855 13970 20919
rect 14034 20855 14858 20919
rect 12300 20825 14858 20855
rect 12300 20761 13281 20825
rect 13345 20761 13371 20825
rect 13435 20761 13461 20825
rect 13525 20761 13551 20825
rect 13615 20761 13640 20825
rect 13704 20823 14858 20825
rect 13704 20761 13749 20823
rect 12300 20759 13749 20761
rect 13813 20816 14858 20823
rect 13813 20759 13851 20816
rect 12300 20752 13851 20759
rect 13915 20752 14858 20816
rect 12300 20712 14858 20752
rect 12300 20709 13749 20712
rect 12300 20645 13281 20709
rect 13345 20645 13371 20709
rect 13435 20645 13461 20709
rect 13525 20645 13551 20709
rect 13615 20645 13640 20709
rect 13704 20648 13749 20709
rect 13813 20648 14858 20712
rect 13704 20645 14858 20648
rect 12300 20631 14858 20645
rect 12300 20567 13140 20631
rect 13204 20593 14858 20631
rect 13204 20567 13281 20593
rect 12300 20529 13281 20567
rect 13345 20529 13371 20593
rect 13435 20529 13461 20593
rect 13525 20529 13551 20593
rect 13615 20529 13640 20593
rect 13704 20529 14858 20593
rect 12300 20505 14858 20529
rect 12300 20441 12961 20505
rect 13025 20441 13051 20505
rect 13115 20441 13141 20505
rect 13205 20441 13231 20505
rect 13295 20441 13320 20505
rect 13384 20469 14858 20505
rect 13384 20441 13428 20469
rect 12300 20405 13428 20441
rect 13492 20405 14858 20469
rect 12300 20389 14858 20405
rect 12300 20325 12961 20389
rect 13025 20325 13051 20389
rect 13115 20325 13141 20389
rect 13205 20325 13231 20389
rect 13295 20325 13320 20389
rect 13384 20325 14858 20389
rect 12300 20306 14858 20325
rect 2055 20209 2700 20242
rect 99 20181 2700 20209
rect 99 20141 1956 20181
rect 99 20077 1852 20141
rect 1916 20117 1956 20141
rect 2020 20117 2045 20181
rect 2109 20117 2135 20181
rect 2199 20117 2225 20181
rect 2289 20117 2315 20181
rect 2379 20117 2700 20181
rect 1916 20077 2700 20117
rect 99 20070 2700 20077
tri 2700 20070 2909 20279 sw
tri 12111 20070 12300 20259 se
rect 12300 20242 12815 20306
rect 12879 20273 14858 20306
rect 12879 20242 12961 20273
rect 12300 20209 12961 20242
rect 13025 20209 13051 20273
rect 13115 20209 13141 20273
rect 13205 20209 13231 20273
rect 13295 20209 13320 20273
rect 13384 20209 14858 20273
rect 12300 20181 14858 20209
rect 12300 20117 12637 20181
rect 12701 20117 12727 20181
rect 12791 20117 12817 20181
rect 12881 20117 12907 20181
rect 12971 20117 12996 20181
rect 13060 20141 14858 20181
rect 13060 20117 13100 20141
rect 12300 20077 13100 20117
rect 13164 20077 14858 20141
rect 12300 20070 14858 20077
rect 99 20065 2456 20070
rect 99 20001 1956 20065
rect 2020 20001 2045 20065
rect 2109 20001 2135 20065
rect 2199 20001 2225 20065
rect 2289 20001 2315 20065
rect 2379 20006 2456 20065
rect 2520 20006 2571 20070
rect 2635 20006 2686 20070
rect 2750 20006 2802 20070
rect 2866 20006 2909 20070
tri 2909 20006 2973 20070 sw
tri 12110 20069 12111 20070 se
rect 12111 20069 12150 20070
tri 12047 20006 12110 20069 se
rect 12110 20006 12150 20069
rect 12214 20006 12266 20070
rect 12330 20006 12381 20070
rect 12445 20006 12496 20070
rect 12560 20065 14858 20070
rect 12560 20006 12637 20065
rect 2379 20001 2973 20006
rect 99 19955 2973 20001
rect 99 19950 2906 19955
rect 99 19949 2456 19950
rect 99 19885 1956 19949
rect 2020 19885 2045 19949
rect 2109 19885 2135 19949
rect 2199 19885 2225 19949
rect 2289 19885 2315 19949
rect 2379 19886 2456 19949
rect 2520 19886 2571 19950
rect 2635 19886 2686 19950
rect 2750 19886 2802 19950
rect 2866 19891 2906 19950
rect 2970 19891 2973 19955
rect 2866 19886 2973 19891
rect 2379 19885 2973 19886
rect 99 19844 2973 19885
tri 2973 19844 3135 20006 sw
tri 12027 19986 12047 20006 se
rect 12047 20001 12637 20006
rect 12701 20001 12727 20065
rect 12791 20001 12817 20065
rect 12881 20001 12907 20065
rect 12971 20001 12996 20065
rect 13060 20001 14858 20065
rect 12047 19986 14858 20001
tri 11885 19844 12027 19986 se
rect 12027 19955 14858 19986
rect 12027 19891 12046 19955
rect 12110 19950 14858 19955
rect 12110 19891 12150 19950
rect 12027 19886 12150 19891
rect 12214 19886 12266 19950
rect 12330 19886 12381 19950
rect 12445 19886 12496 19950
rect 12560 19949 14858 19950
rect 12560 19886 12637 19949
rect 12027 19885 12637 19886
rect 12701 19885 12727 19949
rect 12791 19885 12817 19949
rect 12881 19885 12907 19949
rect 12971 19885 12996 19949
rect 13060 19885 14858 19949
rect 12027 19844 14858 19885
rect 99 19800 2293 19844
rect 99 19736 2193 19800
rect 2257 19780 2293 19800
rect 2357 19780 2377 19844
rect 2441 19780 2461 19844
rect 2525 19780 2545 19844
rect 2609 19780 2629 19844
rect 2693 19780 2713 19844
rect 2777 19780 2797 19844
rect 2861 19780 2881 19844
rect 2945 19780 2965 19844
rect 3029 19780 3049 19844
rect 3113 19780 3135 19844
rect 2257 19736 3135 19780
rect 99 19728 3135 19736
rect 99 19664 2293 19728
rect 2357 19664 2377 19728
rect 2441 19664 2461 19728
rect 2525 19664 2545 19728
rect 2609 19664 2629 19728
rect 2693 19664 2713 19728
rect 2777 19664 2797 19728
rect 2861 19664 2881 19728
rect 2945 19664 2965 19728
rect 3029 19664 3049 19728
rect 3113 19707 3135 19728
tri 3135 19707 3272 19844 sw
tri 11753 19712 11885 19844 se
rect 11885 19780 11903 19844
rect 11967 19780 11987 19844
rect 12051 19780 12071 19844
rect 12135 19780 12155 19844
rect 12219 19780 12239 19844
rect 12303 19780 12323 19844
rect 12387 19780 12407 19844
rect 12471 19780 12491 19844
rect 12555 19780 12575 19844
rect 12639 19780 12659 19844
rect 12723 19800 14858 19844
rect 12723 19780 12759 19800
rect 11885 19736 12759 19780
rect 12823 19736 14858 19800
rect 11885 19728 14858 19736
rect 11885 19712 11903 19728
tri 11748 19707 11753 19712 se
rect 11753 19707 11903 19712
rect 3113 19664 3153 19707
rect 99 19643 3153 19664
rect 3217 19643 3272 19707
rect 99 19614 3272 19643
rect 99 19612 3153 19614
rect 99 19548 2293 19612
rect 2357 19548 2377 19612
rect 2441 19548 2461 19612
rect 2525 19548 2545 19612
rect 2609 19548 2629 19612
rect 2693 19548 2713 19612
rect 2777 19548 2797 19612
rect 2861 19548 2881 19612
rect 2945 19548 2965 19612
rect 3029 19548 3049 19612
rect 3113 19550 3153 19612
rect 3217 19550 3272 19614
rect 3113 19548 3272 19550
rect 99 16575 3272 19548
tri 99 14722 1952 16575 ne
rect 1952 16471 3272 16575
tri 3272 16471 6508 19707 sw
tri 8512 16471 11748 19707 se
rect 11748 19643 11799 19707
rect 11863 19664 11903 19707
rect 11967 19664 11987 19728
rect 12051 19664 12071 19728
rect 12135 19664 12155 19728
rect 12219 19664 12239 19728
rect 12303 19664 12323 19728
rect 12387 19664 12407 19728
rect 12471 19664 12491 19728
rect 12555 19664 12575 19728
rect 12639 19664 12659 19728
rect 12723 19664 14858 19728
rect 11863 19643 14858 19664
rect 11748 19614 14858 19643
rect 11748 19550 11799 19614
rect 11863 19612 14858 19614
rect 11863 19550 11903 19612
rect 11748 19548 11903 19550
rect 11967 19548 11987 19612
rect 12051 19548 12071 19612
rect 12135 19548 12155 19612
rect 12219 19548 12239 19612
rect 12303 19548 12323 19612
rect 12387 19548 12407 19612
rect 12471 19548 12491 19612
rect 12555 19548 12575 19612
rect 12639 19548 12659 19612
rect 12723 19548 14858 19612
rect 11748 16628 14858 19548
rect 11748 16471 12952 16628
rect 1952 14722 12952 16471
tri 12952 14722 14858 16628 nw
tri 1952 11722 4952 14722 ne
rect 4952 11722 9952 14722
tri 9952 11722 12952 14722 nw
rect 3916 10784 5155 10810
rect 3916 10248 3946 10784
rect 5122 10248 5155 10784
rect 858 9756 2098 9787
rect 858 9300 890 9756
rect 2066 9300 2098 9756
rect 858 3611 2098 9300
rect 2396 9501 3635 9528
rect 2396 8965 2427 9501
rect 3603 8965 3635 9501
rect 2396 6025 3635 8965
rect 3916 7963 5155 10248
rect 3916 7419 3977 7963
rect 5081 7419 5155 7963
rect 3916 7345 5155 7419
rect 2396 5241 2423 6025
rect 3607 5241 3635 6025
rect 2396 5122 3635 5241
rect 858 3067 924 3611
rect 2028 3067 2098 3611
rect 858 2999 2098 3067
rect 5552 1 9352 11722
rect 9753 10766 10992 10794
rect 9753 10230 9784 10766
rect 10960 10230 10992 10766
rect 9753 7965 10992 10230
rect 12858 9741 14098 9787
rect 9753 7421 9820 7965
rect 10924 7421 10992 7965
rect 9753 7352 10992 7421
rect 11273 9502 12512 9529
rect 11273 8966 11304 9502
rect 12480 8966 12512 9502
rect 11273 6024 12512 8966
rect 11273 5240 11297 6024
rect 12481 5240 12512 6024
rect 11273 5122 12512 5240
rect 12858 9285 12890 9741
rect 14066 9285 14098 9741
rect 12858 3643 14098 9285
rect 12858 3019 12928 3643
rect 14032 3019 14098 3643
rect 12858 2991 14098 3019
<< via3 >>
rect 2276 34554 2340 34618
rect 2359 34554 2423 34618
rect 2443 34554 2507 34618
rect 2527 34554 2591 34618
rect 2611 34554 2675 34618
rect 2276 34460 2340 34524
rect 2359 34460 2423 34524
rect 2443 34460 2507 34524
rect 2527 34460 2591 34524
rect 2611 34460 2675 34524
rect 2148 34377 2212 34441
rect 2276 34366 2340 34430
rect 2359 34366 2423 34430
rect 2443 34366 2507 34430
rect 2527 34366 2591 34430
rect 2611 34366 2675 34430
rect 2004 34252 2068 34316
rect 2084 34252 2148 34316
rect 2164 34252 2228 34316
rect 2276 34272 2340 34336
rect 2359 34272 2423 34336
rect 2443 34272 2507 34336
rect 2527 34272 2591 34336
rect 2611 34272 2675 34336
rect 1890 34119 1954 34183
rect 2004 34156 2068 34220
rect 2084 34156 2148 34220
rect 2164 34156 2228 34220
rect 2276 34178 2340 34242
rect 2359 34178 2423 34242
rect 2443 34178 2507 34242
rect 2527 34178 2591 34242
rect 2611 34178 2675 34242
rect 2276 34084 2340 34148
rect 2359 34084 2423 34148
rect 2443 34084 2507 34148
rect 2527 34084 2591 34148
rect 2611 34084 2675 34148
rect 1748 34014 1812 34078
rect 1837 34014 1901 34078
rect 1927 34014 1991 34078
rect 2017 34014 2081 34078
rect 2107 34014 2171 34078
rect 1748 33898 1812 33962
rect 1837 33898 1901 33962
rect 1927 33898 1991 33962
rect 2017 33898 2081 33962
rect 2107 33898 2171 33962
rect 2247 33945 2311 34009
rect 1644 33822 1708 33886
rect 1748 33782 1812 33846
rect 1837 33782 1901 33846
rect 1927 33782 1991 33846
rect 2017 33782 2081 33846
rect 2107 33782 2171 33846
rect 1424 33690 1488 33754
rect 1513 33690 1577 33754
rect 1603 33690 1667 33754
rect 1693 33690 1757 33754
rect 1783 33690 1847 33754
rect 1929 33657 1993 33721
rect 1424 33574 1488 33638
rect 1513 33574 1577 33638
rect 1603 33574 1667 33638
rect 1693 33574 1757 33638
rect 1783 33574 1847 33638
rect 1316 33494 1380 33558
rect 1424 33458 1488 33522
rect 1513 33458 1577 33522
rect 1603 33458 1667 33522
rect 1693 33458 1757 33522
rect 1783 33458 1847 33522
rect 12341 34554 12405 34618
rect 12425 34554 12489 34618
rect 12509 34554 12573 34618
rect 12593 34554 12657 34618
rect 12677 34554 12741 34618
rect 12341 34460 12405 34524
rect 12425 34460 12489 34524
rect 12509 34460 12573 34524
rect 12593 34460 12657 34524
rect 12677 34460 12741 34524
rect 12341 34366 12405 34430
rect 12425 34366 12489 34430
rect 12509 34366 12573 34430
rect 12593 34366 12657 34430
rect 12677 34366 12741 34430
rect 12804 34377 12868 34441
rect 12341 34272 12405 34336
rect 12425 34272 12489 34336
rect 12509 34272 12573 34336
rect 12593 34272 12657 34336
rect 12677 34272 12741 34336
rect 12788 34252 12852 34316
rect 12868 34252 12932 34316
rect 12948 34252 13012 34316
rect 12341 34178 12405 34242
rect 12425 34178 12489 34242
rect 12509 34178 12573 34242
rect 12593 34178 12657 34242
rect 12677 34178 12741 34242
rect 12788 34156 12852 34220
rect 12868 34156 12932 34220
rect 12948 34156 13012 34220
rect 12341 34084 12405 34148
rect 12425 34084 12489 34148
rect 12509 34084 12573 34148
rect 12593 34084 12657 34148
rect 12677 34084 12741 34148
rect 13062 34119 13126 34183
rect 12845 34014 12909 34078
rect 12935 34014 12999 34078
rect 13025 34014 13089 34078
rect 13115 34014 13179 34078
rect 13204 34014 13268 34078
rect 12705 33945 12769 34009
rect 12845 33898 12909 33962
rect 12935 33898 12999 33962
rect 13025 33898 13089 33962
rect 13115 33898 13179 33962
rect 13204 33898 13268 33962
rect 12845 33782 12909 33846
rect 12935 33782 12999 33846
rect 13025 33782 13089 33846
rect 13115 33782 13179 33846
rect 13204 33782 13268 33846
rect 13308 33822 13372 33886
rect 13023 33657 13087 33721
rect 13169 33690 13233 33754
rect 13259 33690 13323 33754
rect 13349 33690 13413 33754
rect 13439 33690 13503 33754
rect 13528 33690 13592 33754
rect 13169 33574 13233 33638
rect 13259 33574 13323 33638
rect 13349 33574 13413 33638
rect 13439 33574 13503 33638
rect 13528 33574 13592 33638
rect 13169 33458 13233 33522
rect 13259 33458 13323 33522
rect 13349 33458 13413 33522
rect 13439 33458 13503 33522
rect 13528 33458 13592 33522
rect 13636 33494 13700 33558
rect 1104 33370 1168 33434
rect 1193 33370 1257 33434
rect 1283 33370 1347 33434
rect 1373 33370 1437 33434
rect 1463 33370 1527 33434
rect 1604 33332 1668 33396
rect 1104 33254 1168 33318
rect 1193 33254 1257 33318
rect 1283 33254 1347 33318
rect 1373 33254 1437 33318
rect 1463 33254 1527 33318
rect 1104 33138 1168 33202
rect 1193 33138 1257 33202
rect 1283 33138 1347 33202
rect 1373 33138 1437 33202
rect 1463 33138 1527 33202
rect 982 33045 1046 33109
rect 1072 33045 1136 33109
rect 1162 33045 1226 33109
rect 1252 33045 1316 33109
rect 1342 33045 1406 33109
rect 1432 33045 1496 33109
rect 982 32965 1046 33029
rect 1072 32965 1136 33029
rect 1162 32965 1226 33029
rect 1252 32965 1316 33029
rect 1342 32965 1406 33029
rect 1432 32965 1496 33029
rect 982 32885 1046 32949
rect 1072 32885 1136 32949
rect 1162 32885 1226 32949
rect 1252 32885 1316 32949
rect 1342 32885 1406 32949
rect 1432 32885 1496 32949
rect 982 32805 1046 32869
rect 1072 32805 1136 32869
rect 1162 32805 1226 32869
rect 1252 32805 1316 32869
rect 1342 32805 1406 32869
rect 1432 32805 1496 32869
rect 982 32725 1046 32789
rect 1072 32725 1136 32789
rect 1162 32725 1226 32789
rect 1252 32725 1316 32789
rect 1342 32725 1406 32789
rect 1432 32725 1496 32789
rect 982 32645 1046 32709
rect 1072 32645 1136 32709
rect 1162 32645 1226 32709
rect 1252 32645 1316 32709
rect 1342 32645 1406 32709
rect 1432 32645 1496 32709
rect 982 32565 1046 32629
rect 1072 32565 1136 32629
rect 1162 32565 1226 32629
rect 1252 32565 1316 32629
rect 1342 32565 1406 32629
rect 1432 32565 1496 32629
rect 982 32485 1046 32549
rect 1072 32485 1136 32549
rect 1162 32485 1226 32549
rect 1252 32485 1316 32549
rect 1342 32485 1406 32549
rect 1432 32485 1496 32549
rect 982 32405 1046 32469
rect 1072 32405 1136 32469
rect 1162 32405 1226 32469
rect 1252 32405 1316 32469
rect 1342 32405 1406 32469
rect 1432 32405 1496 32469
rect 982 32325 1046 32389
rect 1072 32325 1136 32389
rect 1162 32325 1226 32389
rect 1252 32325 1316 32389
rect 1342 32325 1406 32389
rect 1432 32325 1496 32389
rect 982 32245 1046 32309
rect 1072 32245 1136 32309
rect 1162 32245 1226 32309
rect 1252 32245 1316 32309
rect 1342 32245 1406 32309
rect 1432 32245 1496 32309
rect 982 32165 1046 32229
rect 1072 32165 1136 32229
rect 1162 32165 1226 32229
rect 1252 32165 1316 32229
rect 1342 32165 1406 32229
rect 1432 32165 1496 32229
rect 982 32085 1046 32149
rect 1072 32085 1136 32149
rect 1162 32085 1226 32149
rect 1252 32085 1316 32149
rect 1342 32085 1406 32149
rect 1432 32085 1496 32149
rect 982 32005 1046 32069
rect 1072 32005 1136 32069
rect 1162 32005 1226 32069
rect 1252 32005 1316 32069
rect 1342 32005 1406 32069
rect 1432 32005 1496 32069
rect 982 31925 1046 31989
rect 1072 31925 1136 31989
rect 1162 31925 1226 31989
rect 1252 31925 1316 31989
rect 1342 31925 1406 31989
rect 1432 31925 1496 31989
rect 982 31845 1046 31909
rect 1072 31845 1136 31909
rect 1162 31845 1226 31909
rect 1252 31845 1316 31909
rect 1342 31845 1406 31909
rect 1432 31845 1496 31909
rect 982 31765 1046 31829
rect 1072 31765 1136 31829
rect 1162 31765 1226 31829
rect 1252 31765 1316 31829
rect 1342 31765 1406 31829
rect 1432 31765 1496 31829
rect 982 31685 1046 31749
rect 1072 31685 1136 31749
rect 1162 31685 1226 31749
rect 1252 31685 1316 31749
rect 1342 31685 1406 31749
rect 1432 31685 1496 31749
rect 982 31605 1046 31669
rect 1072 31605 1136 31669
rect 1162 31605 1226 31669
rect 1252 31605 1316 31669
rect 1342 31605 1406 31669
rect 1432 31605 1496 31669
rect 982 31525 1046 31589
rect 1072 31525 1136 31589
rect 1162 31525 1226 31589
rect 1252 31525 1316 31589
rect 1342 31525 1406 31589
rect 1432 31525 1496 31589
rect 982 31445 1046 31509
rect 1072 31445 1136 31509
rect 1162 31445 1226 31509
rect 1252 31445 1316 31509
rect 1342 31445 1406 31509
rect 1432 31445 1496 31509
rect 982 31365 1046 31429
rect 1072 31365 1136 31429
rect 1162 31365 1226 31429
rect 1252 31365 1316 31429
rect 1342 31365 1406 31429
rect 1432 31365 1496 31429
rect 982 31285 1046 31349
rect 1072 31285 1136 31349
rect 1162 31285 1226 31349
rect 1252 31285 1316 31349
rect 1342 31285 1406 31349
rect 1432 31285 1496 31349
rect 982 31205 1046 31269
rect 1072 31205 1136 31269
rect 1162 31205 1226 31269
rect 1252 31205 1316 31269
rect 1342 31205 1406 31269
rect 1432 31205 1496 31269
rect 982 31125 1046 31189
rect 1072 31125 1136 31189
rect 1162 31125 1226 31189
rect 1252 31125 1316 31189
rect 1342 31125 1406 31189
rect 1432 31125 1496 31189
rect 982 31045 1046 31109
rect 1072 31045 1136 31109
rect 1162 31045 1226 31109
rect 1252 31045 1316 31109
rect 1342 31045 1406 31109
rect 1432 31045 1496 31109
rect 982 30965 1046 31029
rect 1072 30965 1136 31029
rect 1162 30965 1226 31029
rect 1252 30965 1316 31029
rect 1342 30965 1406 31029
rect 1432 30965 1496 31029
rect 982 30885 1046 30949
rect 1072 30885 1136 30949
rect 1162 30885 1226 30949
rect 1252 30885 1316 30949
rect 1342 30885 1406 30949
rect 1432 30885 1496 30949
rect 982 30805 1046 30869
rect 1072 30805 1136 30869
rect 1162 30805 1226 30869
rect 1252 30805 1316 30869
rect 1342 30805 1406 30869
rect 1432 30805 1496 30869
rect 982 30725 1046 30789
rect 1072 30725 1136 30789
rect 1162 30725 1226 30789
rect 1252 30725 1316 30789
rect 1342 30725 1406 30789
rect 1432 30725 1496 30789
rect 982 30645 1046 30709
rect 1072 30645 1136 30709
rect 1162 30645 1226 30709
rect 1252 30645 1316 30709
rect 1342 30645 1406 30709
rect 1432 30645 1496 30709
rect 982 30565 1046 30629
rect 1072 30565 1136 30629
rect 1162 30565 1226 30629
rect 1252 30565 1316 30629
rect 1342 30565 1406 30629
rect 1432 30565 1496 30629
rect 982 30485 1046 30549
rect 1072 30485 1136 30549
rect 1162 30485 1226 30549
rect 1252 30485 1316 30549
rect 1342 30485 1406 30549
rect 1432 30485 1496 30549
rect 982 30405 1046 30469
rect 1072 30405 1136 30469
rect 1162 30405 1226 30469
rect 1252 30405 1316 30469
rect 1342 30405 1406 30469
rect 1432 30405 1496 30469
rect 982 30325 1046 30389
rect 1072 30325 1136 30389
rect 1162 30325 1226 30389
rect 1252 30325 1316 30389
rect 1342 30325 1406 30389
rect 1432 30325 1496 30389
rect 982 30245 1046 30309
rect 1072 30245 1136 30309
rect 1162 30245 1226 30309
rect 1252 30245 1316 30309
rect 1342 30245 1406 30309
rect 1432 30245 1496 30309
rect 982 30165 1046 30229
rect 1072 30165 1136 30229
rect 1162 30165 1226 30229
rect 1252 30165 1316 30229
rect 1342 30165 1406 30229
rect 1432 30165 1496 30229
rect 982 30085 1046 30149
rect 1072 30085 1136 30149
rect 1162 30085 1226 30149
rect 1252 30085 1316 30149
rect 1342 30085 1406 30149
rect 1432 30085 1496 30149
rect 982 30005 1046 30069
rect 1072 30005 1136 30069
rect 1162 30005 1226 30069
rect 1252 30005 1316 30069
rect 1342 30005 1406 30069
rect 1432 30005 1496 30069
rect 982 29925 1046 29989
rect 1072 29925 1136 29989
rect 1162 29925 1226 29989
rect 1252 29925 1316 29989
rect 1342 29925 1406 29989
rect 1432 29925 1496 29989
rect 982 29845 1046 29909
rect 1072 29845 1136 29909
rect 1162 29845 1226 29909
rect 1252 29845 1316 29909
rect 1342 29845 1406 29909
rect 1432 29845 1496 29909
rect 982 29765 1046 29829
rect 1072 29765 1136 29829
rect 1162 29765 1226 29829
rect 1252 29765 1316 29829
rect 1342 29765 1406 29829
rect 1432 29765 1496 29829
rect 982 29685 1046 29749
rect 1072 29685 1136 29749
rect 1162 29685 1226 29749
rect 1252 29685 1316 29749
rect 1342 29685 1406 29749
rect 1432 29685 1496 29749
rect 982 29605 1046 29669
rect 1072 29605 1136 29669
rect 1162 29605 1226 29669
rect 1252 29605 1316 29669
rect 1342 29605 1406 29669
rect 1432 29605 1496 29669
rect 982 29525 1046 29589
rect 1072 29525 1136 29589
rect 1162 29525 1226 29589
rect 1252 29525 1316 29589
rect 1342 29525 1406 29589
rect 1432 29525 1496 29589
rect 982 29445 1046 29509
rect 1072 29445 1136 29509
rect 1162 29445 1226 29509
rect 1252 29445 1316 29509
rect 1342 29445 1406 29509
rect 1432 29445 1496 29509
rect 982 29365 1046 29429
rect 1072 29365 1136 29429
rect 1162 29365 1226 29429
rect 1252 29365 1316 29429
rect 1342 29365 1406 29429
rect 1432 29365 1496 29429
rect 982 29285 1046 29349
rect 1072 29285 1136 29349
rect 1162 29285 1226 29349
rect 1252 29285 1316 29349
rect 1342 29285 1406 29349
rect 1432 29285 1496 29349
rect 982 29205 1046 29269
rect 1072 29205 1136 29269
rect 1162 29205 1226 29269
rect 1252 29205 1316 29269
rect 1342 29205 1406 29269
rect 1432 29205 1496 29269
rect 982 29125 1046 29189
rect 1072 29125 1136 29189
rect 1162 29125 1226 29189
rect 1252 29125 1316 29189
rect 1342 29125 1406 29189
rect 1432 29125 1496 29189
rect 982 29045 1046 29109
rect 1072 29045 1136 29109
rect 1162 29045 1226 29109
rect 1252 29045 1316 29109
rect 1342 29045 1406 29109
rect 1432 29045 1496 29109
rect 982 28965 1046 29029
rect 1072 28965 1136 29029
rect 1162 28965 1226 29029
rect 1252 28965 1316 29029
rect 1342 28965 1406 29029
rect 1432 28965 1496 29029
rect 982 28885 1046 28949
rect 1072 28885 1136 28949
rect 1162 28885 1226 28949
rect 1252 28885 1316 28949
rect 1342 28885 1406 28949
rect 1432 28885 1496 28949
rect 982 28805 1046 28869
rect 1072 28805 1136 28869
rect 1162 28805 1226 28869
rect 1252 28805 1316 28869
rect 1342 28805 1406 28869
rect 1432 28805 1496 28869
rect 982 28725 1046 28789
rect 1072 28725 1136 28789
rect 1162 28725 1226 28789
rect 1252 28725 1316 28789
rect 1342 28725 1406 28789
rect 1432 28725 1496 28789
rect 982 28645 1046 28709
rect 1072 28645 1136 28709
rect 1162 28645 1226 28709
rect 1252 28645 1316 28709
rect 1342 28645 1406 28709
rect 1432 28645 1496 28709
rect 982 28565 1046 28629
rect 1072 28565 1136 28629
rect 1162 28565 1226 28629
rect 1252 28565 1316 28629
rect 1342 28565 1406 28629
rect 1432 28565 1496 28629
rect 982 28485 1046 28549
rect 1072 28485 1136 28549
rect 1162 28485 1226 28549
rect 1252 28485 1316 28549
rect 1342 28485 1406 28549
rect 1432 28485 1496 28549
rect 982 28405 1046 28469
rect 1072 28405 1136 28469
rect 1162 28405 1226 28469
rect 1252 28405 1316 28469
rect 1342 28405 1406 28469
rect 1432 28405 1496 28469
rect 982 28325 1046 28389
rect 1072 28325 1136 28389
rect 1162 28325 1226 28389
rect 1252 28325 1316 28389
rect 1342 28325 1406 28389
rect 1432 28325 1496 28389
rect 982 28245 1046 28309
rect 1072 28245 1136 28309
rect 1162 28245 1226 28309
rect 1252 28245 1316 28309
rect 1342 28245 1406 28309
rect 1432 28245 1496 28309
rect 982 28165 1046 28229
rect 1072 28165 1136 28229
rect 1162 28165 1226 28229
rect 1252 28165 1316 28229
rect 1342 28165 1406 28229
rect 1432 28165 1496 28229
rect 982 28085 1046 28149
rect 1072 28085 1136 28149
rect 1162 28085 1226 28149
rect 1252 28085 1316 28149
rect 1342 28085 1406 28149
rect 1432 28085 1496 28149
rect 982 28005 1046 28069
rect 1072 28005 1136 28069
rect 1162 28005 1226 28069
rect 1252 28005 1316 28069
rect 1342 28005 1406 28069
rect 1432 28005 1496 28069
rect 982 27925 1046 27989
rect 1072 27925 1136 27989
rect 1162 27925 1226 27989
rect 1252 27925 1316 27989
rect 1342 27925 1406 27989
rect 1432 27925 1496 27989
rect 982 27845 1046 27909
rect 1072 27845 1136 27909
rect 1162 27845 1226 27909
rect 1252 27845 1316 27909
rect 1342 27845 1406 27909
rect 1432 27845 1496 27909
rect 982 27765 1046 27829
rect 1072 27765 1136 27829
rect 1162 27765 1226 27829
rect 1252 27765 1316 27829
rect 1342 27765 1406 27829
rect 1432 27765 1496 27829
rect 982 27685 1046 27749
rect 1072 27685 1136 27749
rect 1162 27685 1226 27749
rect 1252 27685 1316 27749
rect 1342 27685 1406 27749
rect 1432 27685 1496 27749
rect 982 27605 1046 27669
rect 1072 27605 1136 27669
rect 1162 27605 1226 27669
rect 1252 27605 1316 27669
rect 1342 27605 1406 27669
rect 1432 27605 1496 27669
rect 982 27525 1046 27589
rect 1072 27525 1136 27589
rect 1162 27525 1226 27589
rect 1252 27525 1316 27589
rect 1342 27525 1406 27589
rect 1432 27525 1496 27589
rect 982 27445 1046 27509
rect 1072 27445 1136 27509
rect 1162 27445 1226 27509
rect 1252 27445 1316 27509
rect 1342 27445 1406 27509
rect 1432 27445 1496 27509
rect 982 27365 1046 27429
rect 1072 27365 1136 27429
rect 1162 27365 1226 27429
rect 1252 27365 1316 27429
rect 1342 27365 1406 27429
rect 1432 27365 1496 27429
rect 982 27285 1046 27349
rect 1072 27285 1136 27349
rect 1162 27285 1226 27349
rect 1252 27285 1316 27349
rect 1342 27285 1406 27349
rect 1432 27285 1496 27349
rect 982 27205 1046 27269
rect 1072 27205 1136 27269
rect 1162 27205 1226 27269
rect 1252 27205 1316 27269
rect 1342 27205 1406 27269
rect 1432 27205 1496 27269
rect 982 27125 1046 27189
rect 1072 27125 1136 27189
rect 1162 27125 1226 27189
rect 1252 27125 1316 27189
rect 1342 27125 1406 27189
rect 1432 27125 1496 27189
rect 982 27045 1046 27109
rect 1072 27045 1136 27109
rect 1162 27045 1226 27109
rect 1252 27045 1316 27109
rect 1342 27045 1406 27109
rect 1432 27045 1496 27109
rect 982 26965 1046 27029
rect 1072 26965 1136 27029
rect 1162 26965 1226 27029
rect 1252 26965 1316 27029
rect 1342 26965 1406 27029
rect 1432 26965 1496 27029
rect 982 26885 1046 26949
rect 1072 26885 1136 26949
rect 1162 26885 1226 26949
rect 1252 26885 1316 26949
rect 1342 26885 1406 26949
rect 1432 26885 1496 26949
rect 982 26805 1046 26869
rect 1072 26805 1136 26869
rect 1162 26805 1226 26869
rect 1252 26805 1316 26869
rect 1342 26805 1406 26869
rect 1432 26805 1496 26869
rect 982 26725 1046 26789
rect 1072 26725 1136 26789
rect 1162 26725 1226 26789
rect 1252 26725 1316 26789
rect 1342 26725 1406 26789
rect 1432 26725 1496 26789
rect 982 26645 1046 26709
rect 1072 26645 1136 26709
rect 1162 26645 1226 26709
rect 1252 26645 1316 26709
rect 1342 26645 1406 26709
rect 1432 26645 1496 26709
rect 982 26565 1046 26629
rect 1072 26565 1136 26629
rect 1162 26565 1226 26629
rect 1252 26565 1316 26629
rect 1342 26565 1406 26629
rect 1432 26565 1496 26629
rect 982 26485 1046 26549
rect 1072 26485 1136 26549
rect 1162 26485 1226 26549
rect 1252 26485 1316 26549
rect 1342 26485 1406 26549
rect 1432 26485 1496 26549
rect 982 26405 1046 26469
rect 1072 26405 1136 26469
rect 1162 26405 1226 26469
rect 1252 26405 1316 26469
rect 1342 26405 1406 26469
rect 1432 26405 1496 26469
rect 982 26325 1046 26389
rect 1072 26325 1136 26389
rect 1162 26325 1226 26389
rect 1252 26325 1316 26389
rect 1342 26325 1406 26389
rect 1432 26325 1496 26389
rect 982 26245 1046 26309
rect 1072 26245 1136 26309
rect 1162 26245 1226 26309
rect 1252 26245 1316 26309
rect 1342 26245 1406 26309
rect 1432 26245 1496 26309
rect 982 26165 1046 26229
rect 1072 26165 1136 26229
rect 1162 26165 1226 26229
rect 1252 26165 1316 26229
rect 1342 26165 1406 26229
rect 1432 26165 1496 26229
rect 982 26085 1046 26149
rect 1072 26085 1136 26149
rect 1162 26085 1226 26149
rect 1252 26085 1316 26149
rect 1342 26085 1406 26149
rect 1432 26085 1496 26149
rect 982 26005 1046 26069
rect 1072 26005 1136 26069
rect 1162 26005 1226 26069
rect 1252 26005 1316 26069
rect 1342 26005 1406 26069
rect 1432 26005 1496 26069
rect 982 25925 1046 25989
rect 1072 25925 1136 25989
rect 1162 25925 1226 25989
rect 1252 25925 1316 25989
rect 1342 25925 1406 25989
rect 1432 25925 1496 25989
rect 982 25845 1046 25909
rect 1072 25845 1136 25909
rect 1162 25845 1226 25909
rect 1252 25845 1316 25909
rect 1342 25845 1406 25909
rect 1432 25845 1496 25909
rect 982 25765 1046 25829
rect 1072 25765 1136 25829
rect 1162 25765 1226 25829
rect 1252 25765 1316 25829
rect 1342 25765 1406 25829
rect 1432 25765 1496 25829
rect 982 25685 1046 25749
rect 1072 25685 1136 25749
rect 1162 25685 1226 25749
rect 1252 25685 1316 25749
rect 1342 25685 1406 25749
rect 1432 25685 1496 25749
rect 982 25605 1046 25669
rect 1072 25605 1136 25669
rect 1162 25605 1226 25669
rect 1252 25605 1316 25669
rect 1342 25605 1406 25669
rect 1432 25605 1496 25669
rect 982 25525 1046 25589
rect 1072 25525 1136 25589
rect 1162 25525 1226 25589
rect 1252 25525 1316 25589
rect 1342 25525 1406 25589
rect 1432 25525 1496 25589
rect 982 25445 1046 25509
rect 1072 25445 1136 25509
rect 1162 25445 1226 25509
rect 1252 25445 1316 25509
rect 1342 25445 1406 25509
rect 1432 25445 1496 25509
rect 982 25365 1046 25429
rect 1072 25365 1136 25429
rect 1162 25365 1226 25429
rect 1252 25365 1316 25429
rect 1342 25365 1406 25429
rect 1432 25365 1496 25429
rect 982 25285 1046 25349
rect 1072 25285 1136 25349
rect 1162 25285 1226 25349
rect 1252 25285 1316 25349
rect 1342 25285 1406 25349
rect 1432 25285 1496 25349
rect 982 25205 1046 25269
rect 1072 25205 1136 25269
rect 1162 25205 1226 25269
rect 1252 25205 1316 25269
rect 1342 25205 1406 25269
rect 1432 25205 1496 25269
rect 982 25125 1046 25189
rect 1072 25125 1136 25189
rect 1162 25125 1226 25189
rect 1252 25125 1316 25189
rect 1342 25125 1406 25189
rect 1432 25125 1496 25189
rect 982 25045 1046 25109
rect 1072 25045 1136 25109
rect 1162 25045 1226 25109
rect 1252 25045 1316 25109
rect 1342 25045 1406 25109
rect 1432 25045 1496 25109
rect 982 24965 1046 25029
rect 1072 24965 1136 25029
rect 1162 24965 1226 25029
rect 1252 24965 1316 25029
rect 1342 24965 1406 25029
rect 1432 24965 1496 25029
rect 982 24885 1046 24949
rect 1072 24885 1136 24949
rect 1162 24885 1226 24949
rect 1252 24885 1316 24949
rect 1342 24885 1406 24949
rect 1432 24885 1496 24949
rect 982 24805 1046 24869
rect 1072 24805 1136 24869
rect 1162 24805 1226 24869
rect 1252 24805 1316 24869
rect 1342 24805 1406 24869
rect 1432 24805 1496 24869
rect 982 24725 1046 24789
rect 1072 24725 1136 24789
rect 1162 24725 1226 24789
rect 1252 24725 1316 24789
rect 1342 24725 1406 24789
rect 1432 24725 1496 24789
rect 982 24645 1046 24709
rect 1072 24645 1136 24709
rect 1162 24645 1226 24709
rect 1252 24645 1316 24709
rect 1342 24645 1406 24709
rect 1432 24645 1496 24709
rect 982 24565 1046 24629
rect 1072 24565 1136 24629
rect 1162 24565 1226 24629
rect 1252 24565 1316 24629
rect 1342 24565 1406 24629
rect 1432 24565 1496 24629
rect 982 24485 1046 24549
rect 1072 24485 1136 24549
rect 1162 24485 1226 24549
rect 1252 24485 1316 24549
rect 1342 24485 1406 24549
rect 1432 24485 1496 24549
rect 982 24405 1046 24469
rect 1072 24405 1136 24469
rect 1162 24405 1226 24469
rect 1252 24405 1316 24469
rect 1342 24405 1406 24469
rect 1432 24405 1496 24469
rect 982 24325 1046 24389
rect 1072 24325 1136 24389
rect 1162 24325 1226 24389
rect 1252 24325 1316 24389
rect 1342 24325 1406 24389
rect 1432 24325 1496 24389
rect 982 24245 1046 24309
rect 1072 24245 1136 24309
rect 1162 24245 1226 24309
rect 1252 24245 1316 24309
rect 1342 24245 1406 24309
rect 1432 24245 1496 24309
rect 982 24165 1046 24229
rect 1072 24165 1136 24229
rect 1162 24165 1226 24229
rect 1252 24165 1316 24229
rect 1342 24165 1406 24229
rect 1432 24165 1496 24229
rect 982 24085 1046 24149
rect 1072 24085 1136 24149
rect 1162 24085 1226 24149
rect 1252 24085 1316 24149
rect 1342 24085 1406 24149
rect 1432 24085 1496 24149
rect 982 24005 1046 24069
rect 1072 24005 1136 24069
rect 1162 24005 1226 24069
rect 1252 24005 1316 24069
rect 1342 24005 1406 24069
rect 1432 24005 1496 24069
rect 982 23925 1046 23989
rect 1072 23925 1136 23989
rect 1162 23925 1226 23989
rect 1252 23925 1316 23989
rect 1342 23925 1406 23989
rect 1432 23925 1496 23989
rect 982 23845 1046 23909
rect 1072 23845 1136 23909
rect 1162 23845 1226 23909
rect 1252 23845 1316 23909
rect 1342 23845 1406 23909
rect 1432 23845 1496 23909
rect 982 23765 1046 23829
rect 1072 23765 1136 23829
rect 1162 23765 1226 23829
rect 1252 23765 1316 23829
rect 1342 23765 1406 23829
rect 1432 23765 1496 23829
rect 982 23685 1046 23749
rect 1072 23685 1136 23749
rect 1162 23685 1226 23749
rect 1252 23685 1316 23749
rect 1342 23685 1406 23749
rect 1432 23685 1496 23749
rect 982 23605 1046 23669
rect 1072 23605 1136 23669
rect 1162 23605 1226 23669
rect 1252 23605 1316 23669
rect 1342 23605 1406 23669
rect 1432 23605 1496 23669
rect 982 23525 1046 23589
rect 1072 23525 1136 23589
rect 1162 23525 1226 23589
rect 1252 23525 1316 23589
rect 1342 23525 1406 23589
rect 1432 23525 1496 23589
rect 982 23445 1046 23509
rect 1072 23445 1136 23509
rect 1162 23445 1226 23509
rect 1252 23445 1316 23509
rect 1342 23445 1406 23509
rect 1432 23445 1496 23509
rect 982 23365 1046 23429
rect 1072 23365 1136 23429
rect 1162 23365 1226 23429
rect 1252 23365 1316 23429
rect 1342 23365 1406 23429
rect 1432 23365 1496 23429
rect 982 23285 1046 23349
rect 1072 23285 1136 23349
rect 1162 23285 1226 23349
rect 1252 23285 1316 23349
rect 1342 23285 1406 23349
rect 1432 23285 1496 23349
rect 982 23204 1046 23268
rect 1072 23204 1136 23268
rect 1162 23204 1226 23268
rect 1252 23204 1316 23268
rect 1342 23204 1406 23268
rect 1432 23204 1496 23268
rect 982 23123 1046 23187
rect 1072 23123 1136 23187
rect 1162 23123 1226 23187
rect 1252 23123 1316 23187
rect 1342 23123 1406 23187
rect 1432 23123 1496 23187
rect 982 23042 1046 23106
rect 1072 23042 1136 23106
rect 1162 23042 1226 23106
rect 1252 23042 1316 23106
rect 1342 23042 1406 23106
rect 1432 23042 1496 23106
rect 982 22961 1046 23025
rect 1072 22961 1136 23025
rect 1162 22961 1226 23025
rect 1252 22961 1316 23025
rect 1342 22961 1406 23025
rect 1432 22961 1496 23025
rect 982 22880 1046 22944
rect 1072 22880 1136 22944
rect 1162 22880 1226 22944
rect 1252 22880 1316 22944
rect 1342 22880 1406 22944
rect 1432 22880 1496 22944
rect 982 22799 1046 22863
rect 1072 22799 1136 22863
rect 1162 22799 1226 22863
rect 1252 22799 1316 22863
rect 1342 22799 1406 22863
rect 1432 22799 1496 22863
rect 982 22718 1046 22782
rect 1072 22718 1136 22782
rect 1162 22718 1226 22782
rect 1252 22718 1316 22782
rect 1342 22718 1406 22782
rect 1432 22718 1496 22782
rect 982 22637 1046 22701
rect 1072 22637 1136 22701
rect 1162 22637 1226 22701
rect 1252 22637 1316 22701
rect 1342 22637 1406 22701
rect 1432 22637 1496 22701
rect 982 22556 1046 22620
rect 1072 22556 1136 22620
rect 1162 22556 1226 22620
rect 1252 22556 1316 22620
rect 1342 22556 1406 22620
rect 1432 22556 1496 22620
rect 982 22475 1046 22539
rect 1072 22475 1136 22539
rect 1162 22475 1226 22539
rect 1252 22475 1316 22539
rect 1342 22475 1406 22539
rect 1432 22475 1496 22539
rect 982 22394 1046 22458
rect 1072 22394 1136 22458
rect 1162 22394 1226 22458
rect 1252 22394 1316 22458
rect 1342 22394 1406 22458
rect 1432 22394 1496 22458
rect 982 22313 1046 22377
rect 1072 22313 1136 22377
rect 1162 22313 1226 22377
rect 1252 22313 1316 22377
rect 1342 22313 1406 22377
rect 1432 22313 1496 22377
rect 982 22232 1046 22296
rect 1072 22232 1136 22296
rect 1162 22232 1226 22296
rect 1252 22232 1316 22296
rect 1342 22232 1406 22296
rect 1432 22232 1496 22296
rect 982 22151 1046 22215
rect 1072 22151 1136 22215
rect 1162 22151 1226 22215
rect 1252 22151 1316 22215
rect 1342 22151 1406 22215
rect 1432 22151 1496 22215
rect 982 22070 1046 22134
rect 1072 22070 1136 22134
rect 1162 22070 1226 22134
rect 1252 22070 1316 22134
rect 1342 22070 1406 22134
rect 1432 22070 1496 22134
rect 982 21989 1046 22053
rect 1072 21989 1136 22053
rect 1162 21989 1226 22053
rect 1252 21989 1316 22053
rect 1342 21989 1406 22053
rect 1432 21989 1496 22053
rect 982 21908 1046 21972
rect 1072 21908 1136 21972
rect 1162 21908 1226 21972
rect 1252 21908 1316 21972
rect 1342 21908 1406 21972
rect 1432 21908 1496 21972
rect 982 21827 1046 21891
rect 1072 21827 1136 21891
rect 1162 21827 1226 21891
rect 1252 21827 1316 21891
rect 1342 21827 1406 21891
rect 1432 21827 1496 21891
rect 982 21746 1046 21810
rect 1072 21746 1136 21810
rect 1162 21746 1226 21810
rect 1252 21746 1316 21810
rect 1342 21746 1406 21810
rect 1432 21746 1496 21810
rect 982 21665 1046 21729
rect 1072 21665 1136 21729
rect 1162 21665 1226 21729
rect 1252 21665 1316 21729
rect 1342 21665 1406 21729
rect 1432 21665 1496 21729
rect 982 21584 1046 21648
rect 1072 21584 1136 21648
rect 1162 21584 1226 21648
rect 1252 21584 1316 21648
rect 1342 21584 1406 21648
rect 1432 21584 1496 21648
rect 982 21503 1046 21567
rect 1072 21503 1136 21567
rect 1162 21503 1226 21567
rect 1252 21503 1316 21567
rect 1342 21503 1406 21567
rect 1432 21503 1496 21567
rect 982 21422 1046 21486
rect 1072 21422 1136 21486
rect 1162 21422 1226 21486
rect 1252 21422 1316 21486
rect 1342 21422 1406 21486
rect 1432 21422 1496 21486
rect 982 21341 1046 21405
rect 1072 21341 1136 21405
rect 1162 21341 1226 21405
rect 1252 21341 1316 21405
rect 1342 21341 1406 21405
rect 1432 21341 1496 21405
rect 982 21260 1046 21324
rect 1072 21260 1136 21324
rect 1162 21260 1226 21324
rect 1252 21260 1316 21324
rect 1342 21260 1406 21324
rect 1432 21260 1496 21324
rect 982 21179 1046 21243
rect 1072 21179 1136 21243
rect 1162 21179 1226 21243
rect 1252 21179 1316 21243
rect 1342 21179 1406 21243
rect 1432 21179 1496 21243
rect 982 21098 1046 21162
rect 1072 21098 1136 21162
rect 1162 21098 1226 21162
rect 1252 21098 1316 21162
rect 1342 21098 1406 21162
rect 1432 21098 1496 21162
rect 982 21017 1046 21081
rect 1072 21017 1136 21081
rect 1162 21017 1226 21081
rect 1252 21017 1316 21081
rect 1342 21017 1406 21081
rect 1432 21017 1496 21081
rect 982 20936 1046 21000
rect 1072 20936 1136 21000
rect 1162 20936 1226 21000
rect 1252 20936 1316 21000
rect 1342 20936 1406 21000
rect 1432 20936 1496 21000
rect 982 20855 1046 20919
rect 1072 20855 1136 20919
rect 1162 20855 1226 20919
rect 1252 20855 1316 20919
rect 1342 20855 1406 20919
rect 1432 20855 1496 20919
rect 1531 20875 1595 20939
rect 1141 20719 1205 20783
rect 1312 20761 1376 20825
rect 1401 20761 1465 20825
rect 1491 20761 1555 20825
rect 1581 20761 1645 20825
rect 1671 20761 1735 20825
rect 1312 20645 1376 20709
rect 1401 20645 1465 20709
rect 1491 20645 1555 20709
rect 1581 20645 1645 20709
rect 1671 20645 1735 20709
rect 1312 20529 1376 20593
rect 1401 20529 1465 20593
rect 1491 20529 1555 20593
rect 1581 20529 1645 20593
rect 1671 20529 1735 20593
rect 1812 20567 1876 20631
rect 1524 20405 1588 20469
rect 1632 20441 1696 20505
rect 1721 20441 1785 20505
rect 1811 20441 1875 20505
rect 1901 20441 1965 20505
rect 1991 20441 2055 20505
rect 1632 20325 1696 20389
rect 1721 20325 1785 20389
rect 1811 20325 1875 20389
rect 1901 20325 1965 20389
rect 1991 20325 2055 20389
rect 1632 20209 1696 20273
rect 1721 20209 1785 20273
rect 1811 20209 1875 20273
rect 1901 20209 1965 20273
rect 1991 20209 2055 20273
rect 2137 20242 2201 20306
rect 13348 33332 13412 33396
rect 13489 33370 13553 33434
rect 13579 33370 13643 33434
rect 13669 33370 13733 33434
rect 13759 33370 13823 33434
rect 13848 33370 13912 33434
rect 13489 33254 13553 33318
rect 13579 33254 13643 33318
rect 13669 33254 13733 33318
rect 13759 33254 13823 33318
rect 13848 33254 13912 33318
rect 13489 33138 13553 33202
rect 13579 33138 13643 33202
rect 13669 33138 13733 33202
rect 13759 33138 13823 33202
rect 13848 33138 13912 33202
rect 13520 33045 13584 33109
rect 13610 33045 13674 33109
rect 13700 33045 13764 33109
rect 13790 33045 13854 33109
rect 13880 33045 13944 33109
rect 13970 33045 14034 33109
rect 13520 32965 13584 33029
rect 13610 32965 13674 33029
rect 13700 32965 13764 33029
rect 13790 32965 13854 33029
rect 13880 32965 13944 33029
rect 13970 32965 14034 33029
rect 13520 32885 13584 32949
rect 13610 32885 13674 32949
rect 13700 32885 13764 32949
rect 13790 32885 13854 32949
rect 13880 32885 13944 32949
rect 13970 32885 14034 32949
rect 13520 32805 13584 32869
rect 13610 32805 13674 32869
rect 13700 32805 13764 32869
rect 13790 32805 13854 32869
rect 13880 32805 13944 32869
rect 13970 32805 14034 32869
rect 13520 32725 13584 32789
rect 13610 32725 13674 32789
rect 13700 32725 13764 32789
rect 13790 32725 13854 32789
rect 13880 32725 13944 32789
rect 13970 32725 14034 32789
rect 13520 32645 13584 32709
rect 13610 32645 13674 32709
rect 13700 32645 13764 32709
rect 13790 32645 13854 32709
rect 13880 32645 13944 32709
rect 13970 32645 14034 32709
rect 13520 32565 13584 32629
rect 13610 32565 13674 32629
rect 13700 32565 13764 32629
rect 13790 32565 13854 32629
rect 13880 32565 13944 32629
rect 13970 32565 14034 32629
rect 13520 32485 13584 32549
rect 13610 32485 13674 32549
rect 13700 32485 13764 32549
rect 13790 32485 13854 32549
rect 13880 32485 13944 32549
rect 13970 32485 14034 32549
rect 13520 32405 13584 32469
rect 13610 32405 13674 32469
rect 13700 32405 13764 32469
rect 13790 32405 13854 32469
rect 13880 32405 13944 32469
rect 13970 32405 14034 32469
rect 13520 32325 13584 32389
rect 13610 32325 13674 32389
rect 13700 32325 13764 32389
rect 13790 32325 13854 32389
rect 13880 32325 13944 32389
rect 13970 32325 14034 32389
rect 13520 32245 13584 32309
rect 13610 32245 13674 32309
rect 13700 32245 13764 32309
rect 13790 32245 13854 32309
rect 13880 32245 13944 32309
rect 13970 32245 14034 32309
rect 13520 32165 13584 32229
rect 13610 32165 13674 32229
rect 13700 32165 13764 32229
rect 13790 32165 13854 32229
rect 13880 32165 13944 32229
rect 13970 32165 14034 32229
rect 13520 32085 13584 32149
rect 13610 32085 13674 32149
rect 13700 32085 13764 32149
rect 13790 32085 13854 32149
rect 13880 32085 13944 32149
rect 13970 32085 14034 32149
rect 13520 32005 13584 32069
rect 13610 32005 13674 32069
rect 13700 32005 13764 32069
rect 13790 32005 13854 32069
rect 13880 32005 13944 32069
rect 13970 32005 14034 32069
rect 13520 31925 13584 31989
rect 13610 31925 13674 31989
rect 13700 31925 13764 31989
rect 13790 31925 13854 31989
rect 13880 31925 13944 31989
rect 13970 31925 14034 31989
rect 13520 31845 13584 31909
rect 13610 31845 13674 31909
rect 13700 31845 13764 31909
rect 13790 31845 13854 31909
rect 13880 31845 13944 31909
rect 13970 31845 14034 31909
rect 13520 31765 13584 31829
rect 13610 31765 13674 31829
rect 13700 31765 13764 31829
rect 13790 31765 13854 31829
rect 13880 31765 13944 31829
rect 13970 31765 14034 31829
rect 13520 31685 13584 31749
rect 13610 31685 13674 31749
rect 13700 31685 13764 31749
rect 13790 31685 13854 31749
rect 13880 31685 13944 31749
rect 13970 31685 14034 31749
rect 13520 31605 13584 31669
rect 13610 31605 13674 31669
rect 13700 31605 13764 31669
rect 13790 31605 13854 31669
rect 13880 31605 13944 31669
rect 13970 31605 14034 31669
rect 13520 31525 13584 31589
rect 13610 31525 13674 31589
rect 13700 31525 13764 31589
rect 13790 31525 13854 31589
rect 13880 31525 13944 31589
rect 13970 31525 14034 31589
rect 13520 31445 13584 31509
rect 13610 31445 13674 31509
rect 13700 31445 13764 31509
rect 13790 31445 13854 31509
rect 13880 31445 13944 31509
rect 13970 31445 14034 31509
rect 13520 31365 13584 31429
rect 13610 31365 13674 31429
rect 13700 31365 13764 31429
rect 13790 31365 13854 31429
rect 13880 31365 13944 31429
rect 13970 31365 14034 31429
rect 13520 31285 13584 31349
rect 13610 31285 13674 31349
rect 13700 31285 13764 31349
rect 13790 31285 13854 31349
rect 13880 31285 13944 31349
rect 13970 31285 14034 31349
rect 13520 31205 13584 31269
rect 13610 31205 13674 31269
rect 13700 31205 13764 31269
rect 13790 31205 13854 31269
rect 13880 31205 13944 31269
rect 13970 31205 14034 31269
rect 13520 31125 13584 31189
rect 13610 31125 13674 31189
rect 13700 31125 13764 31189
rect 13790 31125 13854 31189
rect 13880 31125 13944 31189
rect 13970 31125 14034 31189
rect 13520 31045 13584 31109
rect 13610 31045 13674 31109
rect 13700 31045 13764 31109
rect 13790 31045 13854 31109
rect 13880 31045 13944 31109
rect 13970 31045 14034 31109
rect 13520 30965 13584 31029
rect 13610 30965 13674 31029
rect 13700 30965 13764 31029
rect 13790 30965 13854 31029
rect 13880 30965 13944 31029
rect 13970 30965 14034 31029
rect 13520 30885 13584 30949
rect 13610 30885 13674 30949
rect 13700 30885 13764 30949
rect 13790 30885 13854 30949
rect 13880 30885 13944 30949
rect 13970 30885 14034 30949
rect 13520 30805 13584 30869
rect 13610 30805 13674 30869
rect 13700 30805 13764 30869
rect 13790 30805 13854 30869
rect 13880 30805 13944 30869
rect 13970 30805 14034 30869
rect 13520 30725 13584 30789
rect 13610 30725 13674 30789
rect 13700 30725 13764 30789
rect 13790 30725 13854 30789
rect 13880 30725 13944 30789
rect 13970 30725 14034 30789
rect 13520 30645 13584 30709
rect 13610 30645 13674 30709
rect 13700 30645 13764 30709
rect 13790 30645 13854 30709
rect 13880 30645 13944 30709
rect 13970 30645 14034 30709
rect 13520 30565 13584 30629
rect 13610 30565 13674 30629
rect 13700 30565 13764 30629
rect 13790 30565 13854 30629
rect 13880 30565 13944 30629
rect 13970 30565 14034 30629
rect 13520 30485 13584 30549
rect 13610 30485 13674 30549
rect 13700 30485 13764 30549
rect 13790 30485 13854 30549
rect 13880 30485 13944 30549
rect 13970 30485 14034 30549
rect 13520 30405 13584 30469
rect 13610 30405 13674 30469
rect 13700 30405 13764 30469
rect 13790 30405 13854 30469
rect 13880 30405 13944 30469
rect 13970 30405 14034 30469
rect 13520 30325 13584 30389
rect 13610 30325 13674 30389
rect 13700 30325 13764 30389
rect 13790 30325 13854 30389
rect 13880 30325 13944 30389
rect 13970 30325 14034 30389
rect 13520 30245 13584 30309
rect 13610 30245 13674 30309
rect 13700 30245 13764 30309
rect 13790 30245 13854 30309
rect 13880 30245 13944 30309
rect 13970 30245 14034 30309
rect 13520 30165 13584 30229
rect 13610 30165 13674 30229
rect 13700 30165 13764 30229
rect 13790 30165 13854 30229
rect 13880 30165 13944 30229
rect 13970 30165 14034 30229
rect 13520 30085 13584 30149
rect 13610 30085 13674 30149
rect 13700 30085 13764 30149
rect 13790 30085 13854 30149
rect 13880 30085 13944 30149
rect 13970 30085 14034 30149
rect 13520 30005 13584 30069
rect 13610 30005 13674 30069
rect 13700 30005 13764 30069
rect 13790 30005 13854 30069
rect 13880 30005 13944 30069
rect 13970 30005 14034 30069
rect 13520 29925 13584 29989
rect 13610 29925 13674 29989
rect 13700 29925 13764 29989
rect 13790 29925 13854 29989
rect 13880 29925 13944 29989
rect 13970 29925 14034 29989
rect 13520 29845 13584 29909
rect 13610 29845 13674 29909
rect 13700 29845 13764 29909
rect 13790 29845 13854 29909
rect 13880 29845 13944 29909
rect 13970 29845 14034 29909
rect 13520 29765 13584 29829
rect 13610 29765 13674 29829
rect 13700 29765 13764 29829
rect 13790 29765 13854 29829
rect 13880 29765 13944 29829
rect 13970 29765 14034 29829
rect 13520 29685 13584 29749
rect 13610 29685 13674 29749
rect 13700 29685 13764 29749
rect 13790 29685 13854 29749
rect 13880 29685 13944 29749
rect 13970 29685 14034 29749
rect 13520 29605 13584 29669
rect 13610 29605 13674 29669
rect 13700 29605 13764 29669
rect 13790 29605 13854 29669
rect 13880 29605 13944 29669
rect 13970 29605 14034 29669
rect 13520 29525 13584 29589
rect 13610 29525 13674 29589
rect 13700 29525 13764 29589
rect 13790 29525 13854 29589
rect 13880 29525 13944 29589
rect 13970 29525 14034 29589
rect 13520 29445 13584 29509
rect 13610 29445 13674 29509
rect 13700 29445 13764 29509
rect 13790 29445 13854 29509
rect 13880 29445 13944 29509
rect 13970 29445 14034 29509
rect 13520 29365 13584 29429
rect 13610 29365 13674 29429
rect 13700 29365 13764 29429
rect 13790 29365 13854 29429
rect 13880 29365 13944 29429
rect 13970 29365 14034 29429
rect 13520 29285 13584 29349
rect 13610 29285 13674 29349
rect 13700 29285 13764 29349
rect 13790 29285 13854 29349
rect 13880 29285 13944 29349
rect 13970 29285 14034 29349
rect 13520 29205 13584 29269
rect 13610 29205 13674 29269
rect 13700 29205 13764 29269
rect 13790 29205 13854 29269
rect 13880 29205 13944 29269
rect 13970 29205 14034 29269
rect 13520 29125 13584 29189
rect 13610 29125 13674 29189
rect 13700 29125 13764 29189
rect 13790 29125 13854 29189
rect 13880 29125 13944 29189
rect 13970 29125 14034 29189
rect 13520 29045 13584 29109
rect 13610 29045 13674 29109
rect 13700 29045 13764 29109
rect 13790 29045 13854 29109
rect 13880 29045 13944 29109
rect 13970 29045 14034 29109
rect 13520 28965 13584 29029
rect 13610 28965 13674 29029
rect 13700 28965 13764 29029
rect 13790 28965 13854 29029
rect 13880 28965 13944 29029
rect 13970 28965 14034 29029
rect 13520 28885 13584 28949
rect 13610 28885 13674 28949
rect 13700 28885 13764 28949
rect 13790 28885 13854 28949
rect 13880 28885 13944 28949
rect 13970 28885 14034 28949
rect 13520 28805 13584 28869
rect 13610 28805 13674 28869
rect 13700 28805 13764 28869
rect 13790 28805 13854 28869
rect 13880 28805 13944 28869
rect 13970 28805 14034 28869
rect 13520 28725 13584 28789
rect 13610 28725 13674 28789
rect 13700 28725 13764 28789
rect 13790 28725 13854 28789
rect 13880 28725 13944 28789
rect 13970 28725 14034 28789
rect 13520 28645 13584 28709
rect 13610 28645 13674 28709
rect 13700 28645 13764 28709
rect 13790 28645 13854 28709
rect 13880 28645 13944 28709
rect 13970 28645 14034 28709
rect 13520 28565 13584 28629
rect 13610 28565 13674 28629
rect 13700 28565 13764 28629
rect 13790 28565 13854 28629
rect 13880 28565 13944 28629
rect 13970 28565 14034 28629
rect 13520 28485 13584 28549
rect 13610 28485 13674 28549
rect 13700 28485 13764 28549
rect 13790 28485 13854 28549
rect 13880 28485 13944 28549
rect 13970 28485 14034 28549
rect 13520 28405 13584 28469
rect 13610 28405 13674 28469
rect 13700 28405 13764 28469
rect 13790 28405 13854 28469
rect 13880 28405 13944 28469
rect 13970 28405 14034 28469
rect 13520 28325 13584 28389
rect 13610 28325 13674 28389
rect 13700 28325 13764 28389
rect 13790 28325 13854 28389
rect 13880 28325 13944 28389
rect 13970 28325 14034 28389
rect 13520 28245 13584 28309
rect 13610 28245 13674 28309
rect 13700 28245 13764 28309
rect 13790 28245 13854 28309
rect 13880 28245 13944 28309
rect 13970 28245 14034 28309
rect 13520 28165 13584 28229
rect 13610 28165 13674 28229
rect 13700 28165 13764 28229
rect 13790 28165 13854 28229
rect 13880 28165 13944 28229
rect 13970 28165 14034 28229
rect 13520 28085 13584 28149
rect 13610 28085 13674 28149
rect 13700 28085 13764 28149
rect 13790 28085 13854 28149
rect 13880 28085 13944 28149
rect 13970 28085 14034 28149
rect 13520 28005 13584 28069
rect 13610 28005 13674 28069
rect 13700 28005 13764 28069
rect 13790 28005 13854 28069
rect 13880 28005 13944 28069
rect 13970 28005 14034 28069
rect 13520 27925 13584 27989
rect 13610 27925 13674 27989
rect 13700 27925 13764 27989
rect 13790 27925 13854 27989
rect 13880 27925 13944 27989
rect 13970 27925 14034 27989
rect 13520 27845 13584 27909
rect 13610 27845 13674 27909
rect 13700 27845 13764 27909
rect 13790 27845 13854 27909
rect 13880 27845 13944 27909
rect 13970 27845 14034 27909
rect 13520 27765 13584 27829
rect 13610 27765 13674 27829
rect 13700 27765 13764 27829
rect 13790 27765 13854 27829
rect 13880 27765 13944 27829
rect 13970 27765 14034 27829
rect 13520 27685 13584 27749
rect 13610 27685 13674 27749
rect 13700 27685 13764 27749
rect 13790 27685 13854 27749
rect 13880 27685 13944 27749
rect 13970 27685 14034 27749
rect 13520 27605 13584 27669
rect 13610 27605 13674 27669
rect 13700 27605 13764 27669
rect 13790 27605 13854 27669
rect 13880 27605 13944 27669
rect 13970 27605 14034 27669
rect 13520 27525 13584 27589
rect 13610 27525 13674 27589
rect 13700 27525 13764 27589
rect 13790 27525 13854 27589
rect 13880 27525 13944 27589
rect 13970 27525 14034 27589
rect 13520 27445 13584 27509
rect 13610 27445 13674 27509
rect 13700 27445 13764 27509
rect 13790 27445 13854 27509
rect 13880 27445 13944 27509
rect 13970 27445 14034 27509
rect 13520 27365 13584 27429
rect 13610 27365 13674 27429
rect 13700 27365 13764 27429
rect 13790 27365 13854 27429
rect 13880 27365 13944 27429
rect 13970 27365 14034 27429
rect 13520 27285 13584 27349
rect 13610 27285 13674 27349
rect 13700 27285 13764 27349
rect 13790 27285 13854 27349
rect 13880 27285 13944 27349
rect 13970 27285 14034 27349
rect 13520 27205 13584 27269
rect 13610 27205 13674 27269
rect 13700 27205 13764 27269
rect 13790 27205 13854 27269
rect 13880 27205 13944 27269
rect 13970 27205 14034 27269
rect 13520 27125 13584 27189
rect 13610 27125 13674 27189
rect 13700 27125 13764 27189
rect 13790 27125 13854 27189
rect 13880 27125 13944 27189
rect 13970 27125 14034 27189
rect 13520 27045 13584 27109
rect 13610 27045 13674 27109
rect 13700 27045 13764 27109
rect 13790 27045 13854 27109
rect 13880 27045 13944 27109
rect 13970 27045 14034 27109
rect 13520 26965 13584 27029
rect 13610 26965 13674 27029
rect 13700 26965 13764 27029
rect 13790 26965 13854 27029
rect 13880 26965 13944 27029
rect 13970 26965 14034 27029
rect 13520 26885 13584 26949
rect 13610 26885 13674 26949
rect 13700 26885 13764 26949
rect 13790 26885 13854 26949
rect 13880 26885 13944 26949
rect 13970 26885 14034 26949
rect 13520 26805 13584 26869
rect 13610 26805 13674 26869
rect 13700 26805 13764 26869
rect 13790 26805 13854 26869
rect 13880 26805 13944 26869
rect 13970 26805 14034 26869
rect 13520 26725 13584 26789
rect 13610 26725 13674 26789
rect 13700 26725 13764 26789
rect 13790 26725 13854 26789
rect 13880 26725 13944 26789
rect 13970 26725 14034 26789
rect 13520 26645 13584 26709
rect 13610 26645 13674 26709
rect 13700 26645 13764 26709
rect 13790 26645 13854 26709
rect 13880 26645 13944 26709
rect 13970 26645 14034 26709
rect 13520 26565 13584 26629
rect 13610 26565 13674 26629
rect 13700 26565 13764 26629
rect 13790 26565 13854 26629
rect 13880 26565 13944 26629
rect 13970 26565 14034 26629
rect 13520 26485 13584 26549
rect 13610 26485 13674 26549
rect 13700 26485 13764 26549
rect 13790 26485 13854 26549
rect 13880 26485 13944 26549
rect 13970 26485 14034 26549
rect 13520 26405 13584 26469
rect 13610 26405 13674 26469
rect 13700 26405 13764 26469
rect 13790 26405 13854 26469
rect 13880 26405 13944 26469
rect 13970 26405 14034 26469
rect 13520 26325 13584 26389
rect 13610 26325 13674 26389
rect 13700 26325 13764 26389
rect 13790 26325 13854 26389
rect 13880 26325 13944 26389
rect 13970 26325 14034 26389
rect 13520 26245 13584 26309
rect 13610 26245 13674 26309
rect 13700 26245 13764 26309
rect 13790 26245 13854 26309
rect 13880 26245 13944 26309
rect 13970 26245 14034 26309
rect 13520 26165 13584 26229
rect 13610 26165 13674 26229
rect 13700 26165 13764 26229
rect 13790 26165 13854 26229
rect 13880 26165 13944 26229
rect 13970 26165 14034 26229
rect 13520 26085 13584 26149
rect 13610 26085 13674 26149
rect 13700 26085 13764 26149
rect 13790 26085 13854 26149
rect 13880 26085 13944 26149
rect 13970 26085 14034 26149
rect 13520 26005 13584 26069
rect 13610 26005 13674 26069
rect 13700 26005 13764 26069
rect 13790 26005 13854 26069
rect 13880 26005 13944 26069
rect 13970 26005 14034 26069
rect 13520 25925 13584 25989
rect 13610 25925 13674 25989
rect 13700 25925 13764 25989
rect 13790 25925 13854 25989
rect 13880 25925 13944 25989
rect 13970 25925 14034 25989
rect 13520 25845 13584 25909
rect 13610 25845 13674 25909
rect 13700 25845 13764 25909
rect 13790 25845 13854 25909
rect 13880 25845 13944 25909
rect 13970 25845 14034 25909
rect 13520 25765 13584 25829
rect 13610 25765 13674 25829
rect 13700 25765 13764 25829
rect 13790 25765 13854 25829
rect 13880 25765 13944 25829
rect 13970 25765 14034 25829
rect 13520 25685 13584 25749
rect 13610 25685 13674 25749
rect 13700 25685 13764 25749
rect 13790 25685 13854 25749
rect 13880 25685 13944 25749
rect 13970 25685 14034 25749
rect 13520 25605 13584 25669
rect 13610 25605 13674 25669
rect 13700 25605 13764 25669
rect 13790 25605 13854 25669
rect 13880 25605 13944 25669
rect 13970 25605 14034 25669
rect 13520 25525 13584 25589
rect 13610 25525 13674 25589
rect 13700 25525 13764 25589
rect 13790 25525 13854 25589
rect 13880 25525 13944 25589
rect 13970 25525 14034 25589
rect 13520 25445 13584 25509
rect 13610 25445 13674 25509
rect 13700 25445 13764 25509
rect 13790 25445 13854 25509
rect 13880 25445 13944 25509
rect 13970 25445 14034 25509
rect 13520 25365 13584 25429
rect 13610 25365 13674 25429
rect 13700 25365 13764 25429
rect 13790 25365 13854 25429
rect 13880 25365 13944 25429
rect 13970 25365 14034 25429
rect 13520 25285 13584 25349
rect 13610 25285 13674 25349
rect 13700 25285 13764 25349
rect 13790 25285 13854 25349
rect 13880 25285 13944 25349
rect 13970 25285 14034 25349
rect 13520 25205 13584 25269
rect 13610 25205 13674 25269
rect 13700 25205 13764 25269
rect 13790 25205 13854 25269
rect 13880 25205 13944 25269
rect 13970 25205 14034 25269
rect 13520 25125 13584 25189
rect 13610 25125 13674 25189
rect 13700 25125 13764 25189
rect 13790 25125 13854 25189
rect 13880 25125 13944 25189
rect 13970 25125 14034 25189
rect 13520 25045 13584 25109
rect 13610 25045 13674 25109
rect 13700 25045 13764 25109
rect 13790 25045 13854 25109
rect 13880 25045 13944 25109
rect 13970 25045 14034 25109
rect 13520 24965 13584 25029
rect 13610 24965 13674 25029
rect 13700 24965 13764 25029
rect 13790 24965 13854 25029
rect 13880 24965 13944 25029
rect 13970 24965 14034 25029
rect 13520 24885 13584 24949
rect 13610 24885 13674 24949
rect 13700 24885 13764 24949
rect 13790 24885 13854 24949
rect 13880 24885 13944 24949
rect 13970 24885 14034 24949
rect 13520 24805 13584 24869
rect 13610 24805 13674 24869
rect 13700 24805 13764 24869
rect 13790 24805 13854 24869
rect 13880 24805 13944 24869
rect 13970 24805 14034 24869
rect 13520 24725 13584 24789
rect 13610 24725 13674 24789
rect 13700 24725 13764 24789
rect 13790 24725 13854 24789
rect 13880 24725 13944 24789
rect 13970 24725 14034 24789
rect 13520 24645 13584 24709
rect 13610 24645 13674 24709
rect 13700 24645 13764 24709
rect 13790 24645 13854 24709
rect 13880 24645 13944 24709
rect 13970 24645 14034 24709
rect 13520 24565 13584 24629
rect 13610 24565 13674 24629
rect 13700 24565 13764 24629
rect 13790 24565 13854 24629
rect 13880 24565 13944 24629
rect 13970 24565 14034 24629
rect 13520 24485 13584 24549
rect 13610 24485 13674 24549
rect 13700 24485 13764 24549
rect 13790 24485 13854 24549
rect 13880 24485 13944 24549
rect 13970 24485 14034 24549
rect 13520 24405 13584 24469
rect 13610 24405 13674 24469
rect 13700 24405 13764 24469
rect 13790 24405 13854 24469
rect 13880 24405 13944 24469
rect 13970 24405 14034 24469
rect 13520 24325 13584 24389
rect 13610 24325 13674 24389
rect 13700 24325 13764 24389
rect 13790 24325 13854 24389
rect 13880 24325 13944 24389
rect 13970 24325 14034 24389
rect 13520 24245 13584 24309
rect 13610 24245 13674 24309
rect 13700 24245 13764 24309
rect 13790 24245 13854 24309
rect 13880 24245 13944 24309
rect 13970 24245 14034 24309
rect 13520 24165 13584 24229
rect 13610 24165 13674 24229
rect 13700 24165 13764 24229
rect 13790 24165 13854 24229
rect 13880 24165 13944 24229
rect 13970 24165 14034 24229
rect 13520 24085 13584 24149
rect 13610 24085 13674 24149
rect 13700 24085 13764 24149
rect 13790 24085 13854 24149
rect 13880 24085 13944 24149
rect 13970 24085 14034 24149
rect 13520 24005 13584 24069
rect 13610 24005 13674 24069
rect 13700 24005 13764 24069
rect 13790 24005 13854 24069
rect 13880 24005 13944 24069
rect 13970 24005 14034 24069
rect 13520 23925 13584 23989
rect 13610 23925 13674 23989
rect 13700 23925 13764 23989
rect 13790 23925 13854 23989
rect 13880 23925 13944 23989
rect 13970 23925 14034 23989
rect 13520 23845 13584 23909
rect 13610 23845 13674 23909
rect 13700 23845 13764 23909
rect 13790 23845 13854 23909
rect 13880 23845 13944 23909
rect 13970 23845 14034 23909
rect 13520 23765 13584 23829
rect 13610 23765 13674 23829
rect 13700 23765 13764 23829
rect 13790 23765 13854 23829
rect 13880 23765 13944 23829
rect 13970 23765 14034 23829
rect 13520 23685 13584 23749
rect 13610 23685 13674 23749
rect 13700 23685 13764 23749
rect 13790 23685 13854 23749
rect 13880 23685 13944 23749
rect 13970 23685 14034 23749
rect 13520 23605 13584 23669
rect 13610 23605 13674 23669
rect 13700 23605 13764 23669
rect 13790 23605 13854 23669
rect 13880 23605 13944 23669
rect 13970 23605 14034 23669
rect 13520 23525 13584 23589
rect 13610 23525 13674 23589
rect 13700 23525 13764 23589
rect 13790 23525 13854 23589
rect 13880 23525 13944 23589
rect 13970 23525 14034 23589
rect 13520 23445 13584 23509
rect 13610 23445 13674 23509
rect 13700 23445 13764 23509
rect 13790 23445 13854 23509
rect 13880 23445 13944 23509
rect 13970 23445 14034 23509
rect 13520 23365 13584 23429
rect 13610 23365 13674 23429
rect 13700 23365 13764 23429
rect 13790 23365 13854 23429
rect 13880 23365 13944 23429
rect 13970 23365 14034 23429
rect 13520 23285 13584 23349
rect 13610 23285 13674 23349
rect 13700 23285 13764 23349
rect 13790 23285 13854 23349
rect 13880 23285 13944 23349
rect 13970 23285 14034 23349
rect 13520 23204 13584 23268
rect 13610 23204 13674 23268
rect 13700 23204 13764 23268
rect 13790 23204 13854 23268
rect 13880 23204 13944 23268
rect 13970 23204 14034 23268
rect 13520 23123 13584 23187
rect 13610 23123 13674 23187
rect 13700 23123 13764 23187
rect 13790 23123 13854 23187
rect 13880 23123 13944 23187
rect 13970 23123 14034 23187
rect 13520 23042 13584 23106
rect 13610 23042 13674 23106
rect 13700 23042 13764 23106
rect 13790 23042 13854 23106
rect 13880 23042 13944 23106
rect 13970 23042 14034 23106
rect 13520 22961 13584 23025
rect 13610 22961 13674 23025
rect 13700 22961 13764 23025
rect 13790 22961 13854 23025
rect 13880 22961 13944 23025
rect 13970 22961 14034 23025
rect 13520 22880 13584 22944
rect 13610 22880 13674 22944
rect 13700 22880 13764 22944
rect 13790 22880 13854 22944
rect 13880 22880 13944 22944
rect 13970 22880 14034 22944
rect 13520 22799 13584 22863
rect 13610 22799 13674 22863
rect 13700 22799 13764 22863
rect 13790 22799 13854 22863
rect 13880 22799 13944 22863
rect 13970 22799 14034 22863
rect 13520 22718 13584 22782
rect 13610 22718 13674 22782
rect 13700 22718 13764 22782
rect 13790 22718 13854 22782
rect 13880 22718 13944 22782
rect 13970 22718 14034 22782
rect 13520 22637 13584 22701
rect 13610 22637 13674 22701
rect 13700 22637 13764 22701
rect 13790 22637 13854 22701
rect 13880 22637 13944 22701
rect 13970 22637 14034 22701
rect 13520 22556 13584 22620
rect 13610 22556 13674 22620
rect 13700 22556 13764 22620
rect 13790 22556 13854 22620
rect 13880 22556 13944 22620
rect 13970 22556 14034 22620
rect 13520 22475 13584 22539
rect 13610 22475 13674 22539
rect 13700 22475 13764 22539
rect 13790 22475 13854 22539
rect 13880 22475 13944 22539
rect 13970 22475 14034 22539
rect 13520 22394 13584 22458
rect 13610 22394 13674 22458
rect 13700 22394 13764 22458
rect 13790 22394 13854 22458
rect 13880 22394 13944 22458
rect 13970 22394 14034 22458
rect 13520 22313 13584 22377
rect 13610 22313 13674 22377
rect 13700 22313 13764 22377
rect 13790 22313 13854 22377
rect 13880 22313 13944 22377
rect 13970 22313 14034 22377
rect 13520 22232 13584 22296
rect 13610 22232 13674 22296
rect 13700 22232 13764 22296
rect 13790 22232 13854 22296
rect 13880 22232 13944 22296
rect 13970 22232 14034 22296
rect 13520 22151 13584 22215
rect 13610 22151 13674 22215
rect 13700 22151 13764 22215
rect 13790 22151 13854 22215
rect 13880 22151 13944 22215
rect 13970 22151 14034 22215
rect 13520 22070 13584 22134
rect 13610 22070 13674 22134
rect 13700 22070 13764 22134
rect 13790 22070 13854 22134
rect 13880 22070 13944 22134
rect 13970 22070 14034 22134
rect 13520 21989 13584 22053
rect 13610 21989 13674 22053
rect 13700 21989 13764 22053
rect 13790 21989 13854 22053
rect 13880 21989 13944 22053
rect 13970 21989 14034 22053
rect 13520 21908 13584 21972
rect 13610 21908 13674 21972
rect 13700 21908 13764 21972
rect 13790 21908 13854 21972
rect 13880 21908 13944 21972
rect 13970 21908 14034 21972
rect 13520 21827 13584 21891
rect 13610 21827 13674 21891
rect 13700 21827 13764 21891
rect 13790 21827 13854 21891
rect 13880 21827 13944 21891
rect 13970 21827 14034 21891
rect 13520 21746 13584 21810
rect 13610 21746 13674 21810
rect 13700 21746 13764 21810
rect 13790 21746 13854 21810
rect 13880 21746 13944 21810
rect 13970 21746 14034 21810
rect 13520 21665 13584 21729
rect 13610 21665 13674 21729
rect 13700 21665 13764 21729
rect 13790 21665 13854 21729
rect 13880 21665 13944 21729
rect 13970 21665 14034 21729
rect 13520 21584 13584 21648
rect 13610 21584 13674 21648
rect 13700 21584 13764 21648
rect 13790 21584 13854 21648
rect 13880 21584 13944 21648
rect 13970 21584 14034 21648
rect 13520 21503 13584 21567
rect 13610 21503 13674 21567
rect 13700 21503 13764 21567
rect 13790 21503 13854 21567
rect 13880 21503 13944 21567
rect 13970 21503 14034 21567
rect 13520 21422 13584 21486
rect 13610 21422 13674 21486
rect 13700 21422 13764 21486
rect 13790 21422 13854 21486
rect 13880 21422 13944 21486
rect 13970 21422 14034 21486
rect 13520 21341 13584 21405
rect 13610 21341 13674 21405
rect 13700 21341 13764 21405
rect 13790 21341 13854 21405
rect 13880 21341 13944 21405
rect 13970 21341 14034 21405
rect 13520 21260 13584 21324
rect 13610 21260 13674 21324
rect 13700 21260 13764 21324
rect 13790 21260 13854 21324
rect 13880 21260 13944 21324
rect 13970 21260 14034 21324
rect 13520 21179 13584 21243
rect 13610 21179 13674 21243
rect 13700 21179 13764 21243
rect 13790 21179 13854 21243
rect 13880 21179 13944 21243
rect 13970 21179 14034 21243
rect 13520 21098 13584 21162
rect 13610 21098 13674 21162
rect 13700 21098 13764 21162
rect 13790 21098 13854 21162
rect 13880 21098 13944 21162
rect 13970 21098 14034 21162
rect 13520 21017 13584 21081
rect 13610 21017 13674 21081
rect 13700 21017 13764 21081
rect 13790 21017 13854 21081
rect 13880 21017 13944 21081
rect 13970 21017 14034 21081
rect 13421 20875 13485 20939
rect 13520 20936 13584 21000
rect 13610 20936 13674 21000
rect 13700 20936 13764 21000
rect 13790 20936 13854 21000
rect 13880 20936 13944 21000
rect 13970 20936 14034 21000
rect 13520 20855 13584 20919
rect 13610 20855 13674 20919
rect 13700 20855 13764 20919
rect 13790 20855 13854 20919
rect 13880 20855 13944 20919
rect 13970 20855 14034 20919
rect 13281 20761 13345 20825
rect 13371 20761 13435 20825
rect 13461 20761 13525 20825
rect 13551 20761 13615 20825
rect 13640 20761 13704 20825
rect 13749 20759 13813 20823
rect 13851 20752 13915 20816
rect 13281 20645 13345 20709
rect 13371 20645 13435 20709
rect 13461 20645 13525 20709
rect 13551 20645 13615 20709
rect 13640 20645 13704 20709
rect 13749 20648 13813 20712
rect 13140 20567 13204 20631
rect 13281 20529 13345 20593
rect 13371 20529 13435 20593
rect 13461 20529 13525 20593
rect 13551 20529 13615 20593
rect 13640 20529 13704 20593
rect 12961 20441 13025 20505
rect 13051 20441 13115 20505
rect 13141 20441 13205 20505
rect 13231 20441 13295 20505
rect 13320 20441 13384 20505
rect 13428 20405 13492 20469
rect 12961 20325 13025 20389
rect 13051 20325 13115 20389
rect 13141 20325 13205 20389
rect 13231 20325 13295 20389
rect 13320 20325 13384 20389
rect 1852 20077 1916 20141
rect 1956 20117 2020 20181
rect 2045 20117 2109 20181
rect 2135 20117 2199 20181
rect 2225 20117 2289 20181
rect 2315 20117 2379 20181
rect 12815 20242 12879 20306
rect 12961 20209 13025 20273
rect 13051 20209 13115 20273
rect 13141 20209 13205 20273
rect 13231 20209 13295 20273
rect 13320 20209 13384 20273
rect 12637 20117 12701 20181
rect 12727 20117 12791 20181
rect 12817 20117 12881 20181
rect 12907 20117 12971 20181
rect 12996 20117 13060 20181
rect 13100 20077 13164 20141
rect 1956 20001 2020 20065
rect 2045 20001 2109 20065
rect 2135 20001 2199 20065
rect 2225 20001 2289 20065
rect 2315 20001 2379 20065
rect 2456 20006 2520 20070
rect 2571 20006 2635 20070
rect 2686 20006 2750 20070
rect 2802 20006 2866 20070
rect 12150 20006 12214 20070
rect 12266 20006 12330 20070
rect 12381 20006 12445 20070
rect 12496 20006 12560 20070
rect 1956 19885 2020 19949
rect 2045 19885 2109 19949
rect 2135 19885 2199 19949
rect 2225 19885 2289 19949
rect 2315 19885 2379 19949
rect 2456 19886 2520 19950
rect 2571 19886 2635 19950
rect 2686 19886 2750 19950
rect 2802 19886 2866 19950
rect 2906 19891 2970 19955
rect 12637 20001 12701 20065
rect 12727 20001 12791 20065
rect 12817 20001 12881 20065
rect 12907 20001 12971 20065
rect 12996 20001 13060 20065
rect 12046 19891 12110 19955
rect 12150 19886 12214 19950
rect 12266 19886 12330 19950
rect 12381 19886 12445 19950
rect 12496 19886 12560 19950
rect 12637 19885 12701 19949
rect 12727 19885 12791 19949
rect 12817 19885 12881 19949
rect 12907 19885 12971 19949
rect 12996 19885 13060 19949
rect 2193 19736 2257 19800
rect 2293 19780 2357 19844
rect 2377 19780 2441 19844
rect 2461 19780 2525 19844
rect 2545 19780 2609 19844
rect 2629 19780 2693 19844
rect 2713 19780 2777 19844
rect 2797 19780 2861 19844
rect 2881 19780 2945 19844
rect 2965 19780 3029 19844
rect 3049 19780 3113 19844
rect 2293 19664 2357 19728
rect 2377 19664 2441 19728
rect 2461 19664 2525 19728
rect 2545 19664 2609 19728
rect 2629 19664 2693 19728
rect 2713 19664 2777 19728
rect 2797 19664 2861 19728
rect 2881 19664 2945 19728
rect 2965 19664 3029 19728
rect 3049 19664 3113 19728
rect 11903 19780 11967 19844
rect 11987 19780 12051 19844
rect 12071 19780 12135 19844
rect 12155 19780 12219 19844
rect 12239 19780 12303 19844
rect 12323 19780 12387 19844
rect 12407 19780 12471 19844
rect 12491 19780 12555 19844
rect 12575 19780 12639 19844
rect 12659 19780 12723 19844
rect 12759 19736 12823 19800
rect 3153 19643 3217 19707
rect 2293 19548 2357 19612
rect 2377 19548 2441 19612
rect 2461 19548 2525 19612
rect 2545 19548 2609 19612
rect 2629 19548 2693 19612
rect 2713 19548 2777 19612
rect 2797 19548 2861 19612
rect 2881 19548 2945 19612
rect 2965 19548 3029 19612
rect 3049 19548 3113 19612
rect 3153 19550 3217 19614
rect 11799 19643 11863 19707
rect 11903 19664 11967 19728
rect 11987 19664 12051 19728
rect 12071 19664 12135 19728
rect 12155 19664 12219 19728
rect 12239 19664 12303 19728
rect 12323 19664 12387 19728
rect 12407 19664 12471 19728
rect 12491 19664 12555 19728
rect 12575 19664 12639 19728
rect 12659 19664 12723 19728
rect 11799 19550 11863 19614
rect 11903 19548 11967 19612
rect 11987 19548 12051 19612
rect 12071 19548 12135 19612
rect 12155 19548 12219 19612
rect 12239 19548 12303 19612
rect 12323 19548 12387 19612
rect 12407 19548 12471 19612
rect 12491 19548 12555 19612
rect 12575 19548 12639 19612
rect 12659 19548 12723 19612
rect 3977 7419 5081 7963
rect 2423 5241 3607 6025
rect 924 3067 2028 3611
rect 9820 7421 10924 7965
rect 11297 5240 12481 6024
rect 12928 3019 14032 3643
<< metal4 >>
rect 767 36409 1727 37008
rect 13204 36409 14164 37008
rect 2275 34618 2676 34621
rect 2275 34554 2276 34618
rect 2340 34554 2359 34618
rect 2423 34554 2443 34618
rect 2507 34554 2527 34618
rect 2591 34554 2611 34618
rect 2675 34554 2676 34618
rect 2275 34524 2676 34554
rect 2131 34441 2213 34474
rect 2131 34377 2148 34441
rect 2212 34377 2213 34441
rect 2131 34344 2213 34377
rect 2275 34460 2276 34524
rect 2340 34460 2359 34524
rect 2423 34460 2443 34524
rect 2507 34460 2527 34524
rect 2591 34460 2611 34524
rect 2675 34460 2676 34524
rect 2275 34430 2676 34460
rect 2275 34366 2276 34430
rect 2340 34366 2359 34430
rect 2423 34366 2443 34430
rect 2507 34366 2527 34430
rect 2591 34366 2611 34430
rect 2675 34366 2676 34430
rect 2275 34336 2676 34366
rect 2002 34316 2230 34317
rect 2002 34252 2004 34316
rect 2068 34252 2084 34316
rect 2148 34252 2164 34316
rect 2228 34252 2230 34316
rect 2002 34220 2230 34252
rect 1873 34183 1955 34216
rect 1873 34119 1890 34183
rect 1954 34119 1955 34183
rect 2002 34156 2004 34220
rect 2068 34156 2084 34220
rect 2148 34156 2164 34220
rect 2228 34156 2230 34220
rect 2002 34155 2230 34156
rect 2275 34272 2276 34336
rect 2340 34272 2359 34336
rect 2423 34272 2443 34336
rect 2507 34272 2527 34336
rect 2591 34272 2611 34336
rect 2675 34272 2676 34336
rect 2275 34242 2676 34272
rect 2275 34178 2276 34242
rect 2340 34178 2359 34242
rect 2423 34178 2443 34242
rect 2507 34178 2527 34242
rect 2591 34178 2611 34242
rect 2675 34178 2676 34242
rect 1873 34086 1955 34119
rect 2275 34148 2676 34178
rect 2275 34084 2276 34148
rect 2340 34084 2359 34148
rect 2423 34084 2443 34148
rect 2507 34084 2527 34148
rect 2591 34084 2611 34148
rect 2675 34084 2676 34148
rect 2275 34081 2676 34084
rect 12340 34618 12742 34621
rect 12340 34554 12341 34618
rect 12405 34554 12425 34618
rect 12489 34554 12509 34618
rect 12573 34554 12593 34618
rect 12657 34554 12677 34618
rect 12741 34554 12742 34618
rect 12340 34524 12742 34554
rect 12340 34460 12341 34524
rect 12405 34460 12425 34524
rect 12489 34460 12509 34524
rect 12573 34460 12593 34524
rect 12657 34460 12677 34524
rect 12741 34460 12742 34524
rect 12340 34430 12742 34460
rect 12340 34366 12341 34430
rect 12405 34366 12425 34430
rect 12489 34366 12509 34430
rect 12573 34366 12593 34430
rect 12657 34366 12677 34430
rect 12741 34366 12742 34430
rect 12340 34336 12742 34366
rect 12803 34441 12885 34474
rect 12803 34377 12804 34441
rect 12868 34377 12885 34441
rect 12803 34344 12885 34377
rect 12340 34272 12341 34336
rect 12405 34272 12425 34336
rect 12489 34272 12509 34336
rect 12573 34272 12593 34336
rect 12657 34272 12677 34336
rect 12741 34272 12742 34336
rect 12340 34242 12742 34272
rect 12340 34178 12341 34242
rect 12405 34178 12425 34242
rect 12489 34178 12509 34242
rect 12573 34178 12593 34242
rect 12657 34178 12677 34242
rect 12741 34178 12742 34242
rect 12340 34148 12742 34178
rect 12786 34316 13014 34317
rect 12786 34252 12788 34316
rect 12852 34252 12868 34316
rect 12932 34252 12948 34316
rect 13012 34252 13014 34316
rect 12786 34220 13014 34252
rect 12786 34156 12788 34220
rect 12852 34156 12868 34220
rect 12932 34156 12948 34220
rect 13012 34156 13014 34220
rect 12786 34155 13014 34156
rect 13061 34183 13143 34216
rect 12340 34084 12341 34148
rect 12405 34084 12425 34148
rect 12489 34084 12509 34148
rect 12573 34084 12593 34148
rect 12657 34084 12677 34148
rect 12741 34084 12742 34148
rect 13061 34119 13062 34183
rect 13126 34119 13143 34183
rect 13061 34086 13143 34119
rect 12340 34081 12742 34084
rect 1747 34078 2172 34080
rect 1747 34014 1748 34078
rect 1812 34014 1837 34078
rect 1901 34014 1927 34078
rect 1991 34014 2017 34078
rect 2081 34014 2107 34078
rect 2171 34014 2172 34078
rect 12844 34078 13269 34080
rect 1747 33962 2172 34014
rect 1584 33886 1709 33919
rect 1584 33822 1644 33886
rect 1708 33822 1709 33886
rect 1584 33789 1709 33822
rect 1747 33898 1748 33962
rect 1812 33898 1837 33962
rect 1901 33898 1927 33962
rect 1991 33898 2017 33962
rect 2081 33898 2107 33962
rect 2171 33898 2172 33962
rect 2187 34009 2312 34042
rect 2187 33945 2247 34009
rect 2311 33945 2312 34009
rect 2187 33912 2312 33945
rect 12704 34009 12829 34042
rect 12704 33945 12705 34009
rect 12769 33945 12829 34009
rect 12704 33912 12829 33945
rect 12844 34014 12845 34078
rect 12909 34014 12935 34078
rect 12999 34014 13025 34078
rect 13089 34014 13115 34078
rect 13179 34014 13204 34078
rect 13268 34014 13269 34078
rect 12844 33962 13269 34014
rect 1747 33846 2172 33898
rect 1747 33782 1748 33846
rect 1812 33782 1837 33846
rect 1901 33782 1927 33846
rect 1991 33782 2017 33846
rect 2081 33782 2107 33846
rect 2171 33782 2172 33846
rect 1747 33780 2172 33782
rect 12844 33898 12845 33962
rect 12909 33898 12935 33962
rect 12999 33898 13025 33962
rect 13089 33898 13115 33962
rect 13179 33898 13204 33962
rect 13268 33898 13269 33962
rect 12844 33846 13269 33898
rect 12844 33782 12845 33846
rect 12909 33782 12935 33846
rect 12999 33782 13025 33846
rect 13089 33782 13115 33846
rect 13179 33782 13204 33846
rect 13268 33782 13269 33846
rect 13307 33886 13432 33919
rect 13307 33822 13308 33886
rect 13372 33822 13432 33886
rect 13307 33789 13432 33822
rect 12844 33780 13269 33782
rect 1423 33754 1848 33756
rect 13168 33754 13593 33756
rect 1423 33690 1424 33754
rect 1488 33690 1513 33754
rect 1577 33690 1603 33754
rect 1667 33690 1693 33754
rect 1757 33690 1783 33754
rect 1847 33690 1848 33754
rect 1423 33638 1848 33690
rect 1256 33558 1381 33591
rect 1256 33494 1316 33558
rect 1380 33494 1381 33558
rect 1256 33461 1381 33494
rect 1423 33574 1424 33638
rect 1488 33574 1513 33638
rect 1577 33574 1603 33638
rect 1667 33574 1693 33638
rect 1757 33574 1783 33638
rect 1847 33574 1848 33638
rect 1869 33721 1994 33754
rect 1869 33657 1929 33721
rect 1993 33657 1994 33721
rect 1869 33624 1994 33657
rect 13022 33721 13147 33754
rect 13022 33657 13023 33721
rect 13087 33657 13147 33721
rect 13022 33624 13147 33657
rect 13168 33690 13169 33754
rect 13233 33690 13259 33754
rect 13323 33690 13349 33754
rect 13413 33690 13439 33754
rect 13503 33690 13528 33754
rect 13592 33690 13593 33754
rect 13168 33638 13593 33690
rect 1423 33522 1848 33574
rect 1423 33458 1424 33522
rect 1488 33458 1513 33522
rect 1577 33458 1603 33522
rect 1667 33458 1693 33522
rect 1757 33458 1783 33522
rect 1847 33458 1848 33522
rect 1423 33456 1848 33458
rect 13168 33574 13169 33638
rect 13233 33574 13259 33638
rect 13323 33574 13349 33638
rect 13413 33574 13439 33638
rect 13503 33574 13528 33638
rect 13592 33574 13593 33638
rect 13168 33522 13593 33574
rect 13168 33458 13169 33522
rect 13233 33458 13259 33522
rect 13323 33458 13349 33522
rect 13413 33458 13439 33522
rect 13503 33458 13528 33522
rect 13592 33458 13593 33522
rect 13635 33558 13760 33591
rect 13635 33494 13636 33558
rect 13700 33494 13760 33558
rect 13635 33461 13760 33494
rect 13168 33456 13593 33458
rect 1103 33434 1528 33436
rect 1103 33370 1104 33434
rect 1168 33370 1193 33434
rect 1257 33370 1283 33434
rect 1347 33370 1373 33434
rect 1437 33370 1463 33434
rect 1527 33370 1528 33434
rect 13488 33434 13913 33436
rect 1103 33318 1528 33370
rect 1103 33254 1104 33318
rect 1168 33254 1193 33318
rect 1257 33254 1283 33318
rect 1347 33254 1373 33318
rect 1437 33254 1463 33318
rect 1527 33254 1528 33318
rect 1544 33396 1669 33429
rect 1544 33332 1604 33396
rect 1668 33332 1669 33396
rect 1544 33299 1669 33332
rect 13347 33396 13472 33429
rect 13347 33332 13348 33396
rect 13412 33332 13472 33396
rect 13347 33299 13472 33332
rect 13488 33370 13489 33434
rect 13553 33370 13579 33434
rect 13643 33370 13669 33434
rect 13733 33370 13759 33434
rect 13823 33370 13848 33434
rect 13912 33370 13913 33434
rect 13488 33318 13913 33370
rect 1103 33202 1528 33254
rect 1103 33138 1104 33202
rect 1168 33138 1193 33202
rect 1257 33138 1283 33202
rect 1347 33138 1373 33202
rect 1437 33138 1463 33202
rect 1527 33138 1528 33202
rect 1103 33136 1528 33138
rect 13488 33254 13489 33318
rect 13553 33254 13579 33318
rect 13643 33254 13669 33318
rect 13733 33254 13759 33318
rect 13823 33254 13848 33318
rect 13912 33254 13913 33318
rect 13488 33202 13913 33254
rect 13488 33138 13489 33202
rect 13553 33138 13579 33202
rect 13643 33138 13669 33202
rect 13733 33138 13759 33202
rect 13823 33138 13848 33202
rect 13912 33138 13913 33202
rect 13488 33136 13913 33138
rect 977 33109 1501 33110
rect 977 33045 982 33109
rect 1046 33045 1072 33109
rect 1136 33045 1162 33109
rect 1226 33045 1252 33109
rect 1316 33045 1342 33109
rect 1406 33045 1432 33109
rect 1496 33045 1501 33109
rect 977 33029 1501 33045
rect 977 32965 982 33029
rect 1046 32965 1072 33029
rect 1136 32965 1162 33029
rect 1226 32965 1252 33029
rect 1316 32965 1342 33029
rect 1406 32965 1432 33029
rect 1496 32965 1501 33029
rect 977 32949 1501 32965
rect 977 32885 982 32949
rect 1046 32885 1072 32949
rect 1136 32885 1162 32949
rect 1226 32885 1252 32949
rect 1316 32885 1342 32949
rect 1406 32885 1432 32949
rect 1496 32885 1501 32949
rect 977 32869 1501 32885
rect 977 32805 982 32869
rect 1046 32805 1072 32869
rect 1136 32805 1162 32869
rect 1226 32805 1252 32869
rect 1316 32805 1342 32869
rect 1406 32805 1432 32869
rect 1496 32805 1501 32869
rect 977 32789 1501 32805
rect 977 32725 982 32789
rect 1046 32725 1072 32789
rect 1136 32725 1162 32789
rect 1226 32725 1252 32789
rect 1316 32725 1342 32789
rect 1406 32725 1432 32789
rect 1496 32725 1501 32789
rect 977 32709 1501 32725
rect 977 32645 982 32709
rect 1046 32645 1072 32709
rect 1136 32645 1162 32709
rect 1226 32645 1252 32709
rect 1316 32645 1342 32709
rect 1406 32645 1432 32709
rect 1496 32645 1501 32709
rect 977 32629 1501 32645
rect 977 32565 982 32629
rect 1046 32565 1072 32629
rect 1136 32565 1162 32629
rect 1226 32565 1252 32629
rect 1316 32565 1342 32629
rect 1406 32565 1432 32629
rect 1496 32565 1501 32629
rect 977 32549 1501 32565
rect 977 32485 982 32549
rect 1046 32485 1072 32549
rect 1136 32485 1162 32549
rect 1226 32485 1252 32549
rect 1316 32485 1342 32549
rect 1406 32485 1432 32549
rect 1496 32485 1501 32549
rect 977 32469 1501 32485
rect 977 32405 982 32469
rect 1046 32405 1072 32469
rect 1136 32405 1162 32469
rect 1226 32405 1252 32469
rect 1316 32405 1342 32469
rect 1406 32405 1432 32469
rect 1496 32405 1501 32469
rect 977 32389 1501 32405
rect 977 32325 982 32389
rect 1046 32325 1072 32389
rect 1136 32325 1162 32389
rect 1226 32325 1252 32389
rect 1316 32325 1342 32389
rect 1406 32325 1432 32389
rect 1496 32325 1501 32389
rect 977 32309 1501 32325
rect 977 32245 982 32309
rect 1046 32245 1072 32309
rect 1136 32245 1162 32309
rect 1226 32245 1252 32309
rect 1316 32245 1342 32309
rect 1406 32245 1432 32309
rect 1496 32245 1501 32309
rect 977 32229 1501 32245
rect 977 32165 982 32229
rect 1046 32165 1072 32229
rect 1136 32165 1162 32229
rect 1226 32165 1252 32229
rect 1316 32165 1342 32229
rect 1406 32165 1432 32229
rect 1496 32165 1501 32229
rect 977 32149 1501 32165
rect 977 32085 982 32149
rect 1046 32085 1072 32149
rect 1136 32085 1162 32149
rect 1226 32085 1252 32149
rect 1316 32085 1342 32149
rect 1406 32085 1432 32149
rect 1496 32085 1501 32149
rect 977 32069 1501 32085
rect 977 32005 982 32069
rect 1046 32005 1072 32069
rect 1136 32005 1162 32069
rect 1226 32005 1252 32069
rect 1316 32005 1342 32069
rect 1406 32005 1432 32069
rect 1496 32005 1501 32069
rect 977 31989 1501 32005
rect 977 31925 982 31989
rect 1046 31925 1072 31989
rect 1136 31925 1162 31989
rect 1226 31925 1252 31989
rect 1316 31925 1342 31989
rect 1406 31925 1432 31989
rect 1496 31925 1501 31989
rect 977 31909 1501 31925
rect 977 31845 982 31909
rect 1046 31845 1072 31909
rect 1136 31845 1162 31909
rect 1226 31845 1252 31909
rect 1316 31845 1342 31909
rect 1406 31845 1432 31909
rect 1496 31845 1501 31909
rect 977 31829 1501 31845
rect 977 31765 982 31829
rect 1046 31765 1072 31829
rect 1136 31765 1162 31829
rect 1226 31765 1252 31829
rect 1316 31765 1342 31829
rect 1406 31765 1432 31829
rect 1496 31765 1501 31829
rect 977 31749 1501 31765
rect 977 31685 982 31749
rect 1046 31685 1072 31749
rect 1136 31685 1162 31749
rect 1226 31685 1252 31749
rect 1316 31685 1342 31749
rect 1406 31685 1432 31749
rect 1496 31685 1501 31749
rect 977 31669 1501 31685
rect 977 31605 982 31669
rect 1046 31605 1072 31669
rect 1136 31605 1162 31669
rect 1226 31605 1252 31669
rect 1316 31605 1342 31669
rect 1406 31605 1432 31669
rect 1496 31605 1501 31669
rect 977 31589 1501 31605
rect 977 31525 982 31589
rect 1046 31525 1072 31589
rect 1136 31525 1162 31589
rect 1226 31525 1252 31589
rect 1316 31525 1342 31589
rect 1406 31525 1432 31589
rect 1496 31525 1501 31589
rect 977 31509 1501 31525
rect 977 31445 982 31509
rect 1046 31445 1072 31509
rect 1136 31445 1162 31509
rect 1226 31445 1252 31509
rect 1316 31445 1342 31509
rect 1406 31445 1432 31509
rect 1496 31445 1501 31509
rect 977 31429 1501 31445
rect 977 31365 982 31429
rect 1046 31365 1072 31429
rect 1136 31365 1162 31429
rect 1226 31365 1252 31429
rect 1316 31365 1342 31429
rect 1406 31365 1432 31429
rect 1496 31365 1501 31429
rect 977 31349 1501 31365
rect 977 31285 982 31349
rect 1046 31285 1072 31349
rect 1136 31285 1162 31349
rect 1226 31285 1252 31349
rect 1316 31285 1342 31349
rect 1406 31285 1432 31349
rect 1496 31285 1501 31349
rect 977 31269 1501 31285
rect 977 31205 982 31269
rect 1046 31205 1072 31269
rect 1136 31205 1162 31269
rect 1226 31205 1252 31269
rect 1316 31205 1342 31269
rect 1406 31205 1432 31269
rect 1496 31205 1501 31269
rect 977 31189 1501 31205
rect 977 31125 982 31189
rect 1046 31125 1072 31189
rect 1136 31125 1162 31189
rect 1226 31125 1252 31189
rect 1316 31125 1342 31189
rect 1406 31125 1432 31189
rect 1496 31125 1501 31189
rect 977 31109 1501 31125
rect 977 31045 982 31109
rect 1046 31045 1072 31109
rect 1136 31045 1162 31109
rect 1226 31045 1252 31109
rect 1316 31045 1342 31109
rect 1406 31045 1432 31109
rect 1496 31045 1501 31109
rect 977 31029 1501 31045
rect 977 30965 982 31029
rect 1046 30965 1072 31029
rect 1136 30965 1162 31029
rect 1226 30965 1252 31029
rect 1316 30965 1342 31029
rect 1406 30965 1432 31029
rect 1496 30965 1501 31029
rect 977 30949 1501 30965
rect 977 30885 982 30949
rect 1046 30885 1072 30949
rect 1136 30885 1162 30949
rect 1226 30885 1252 30949
rect 1316 30885 1342 30949
rect 1406 30885 1432 30949
rect 1496 30885 1501 30949
rect 977 30869 1501 30885
rect 977 30805 982 30869
rect 1046 30805 1072 30869
rect 1136 30805 1162 30869
rect 1226 30805 1252 30869
rect 1316 30805 1342 30869
rect 1406 30805 1432 30869
rect 1496 30805 1501 30869
rect 977 30789 1501 30805
rect 977 30725 982 30789
rect 1046 30725 1072 30789
rect 1136 30725 1162 30789
rect 1226 30725 1252 30789
rect 1316 30725 1342 30789
rect 1406 30725 1432 30789
rect 1496 30725 1501 30789
rect 977 30709 1501 30725
rect 977 30645 982 30709
rect 1046 30645 1072 30709
rect 1136 30645 1162 30709
rect 1226 30645 1252 30709
rect 1316 30645 1342 30709
rect 1406 30645 1432 30709
rect 1496 30645 1501 30709
rect 977 30629 1501 30645
rect 977 30565 982 30629
rect 1046 30565 1072 30629
rect 1136 30565 1162 30629
rect 1226 30565 1252 30629
rect 1316 30565 1342 30629
rect 1406 30565 1432 30629
rect 1496 30565 1501 30629
rect 977 30549 1501 30565
rect 977 30485 982 30549
rect 1046 30485 1072 30549
rect 1136 30485 1162 30549
rect 1226 30485 1252 30549
rect 1316 30485 1342 30549
rect 1406 30485 1432 30549
rect 1496 30485 1501 30549
rect 977 30469 1501 30485
rect 977 30405 982 30469
rect 1046 30405 1072 30469
rect 1136 30405 1162 30469
rect 1226 30405 1252 30469
rect 1316 30405 1342 30469
rect 1406 30405 1432 30469
rect 1496 30405 1501 30469
rect 977 30389 1501 30405
rect 977 30325 982 30389
rect 1046 30325 1072 30389
rect 1136 30325 1162 30389
rect 1226 30325 1252 30389
rect 1316 30325 1342 30389
rect 1406 30325 1432 30389
rect 1496 30325 1501 30389
rect 977 30309 1501 30325
rect 977 30245 982 30309
rect 1046 30245 1072 30309
rect 1136 30245 1162 30309
rect 1226 30245 1252 30309
rect 1316 30245 1342 30309
rect 1406 30245 1432 30309
rect 1496 30245 1501 30309
rect 977 30229 1501 30245
rect 977 30165 982 30229
rect 1046 30165 1072 30229
rect 1136 30165 1162 30229
rect 1226 30165 1252 30229
rect 1316 30165 1342 30229
rect 1406 30165 1432 30229
rect 1496 30165 1501 30229
rect 977 30149 1501 30165
rect 977 30085 982 30149
rect 1046 30085 1072 30149
rect 1136 30085 1162 30149
rect 1226 30085 1252 30149
rect 1316 30085 1342 30149
rect 1406 30085 1432 30149
rect 1496 30085 1501 30149
rect 977 30069 1501 30085
rect 977 30005 982 30069
rect 1046 30005 1072 30069
rect 1136 30005 1162 30069
rect 1226 30005 1252 30069
rect 1316 30005 1342 30069
rect 1406 30005 1432 30069
rect 1496 30005 1501 30069
rect 977 29989 1501 30005
rect 977 29925 982 29989
rect 1046 29925 1072 29989
rect 1136 29925 1162 29989
rect 1226 29925 1252 29989
rect 1316 29925 1342 29989
rect 1406 29925 1432 29989
rect 1496 29925 1501 29989
rect 977 29909 1501 29925
rect 977 29845 982 29909
rect 1046 29845 1072 29909
rect 1136 29845 1162 29909
rect 1226 29845 1252 29909
rect 1316 29845 1342 29909
rect 1406 29845 1432 29909
rect 1496 29845 1501 29909
rect 977 29829 1501 29845
rect 977 29765 982 29829
rect 1046 29765 1072 29829
rect 1136 29765 1162 29829
rect 1226 29765 1252 29829
rect 1316 29765 1342 29829
rect 1406 29765 1432 29829
rect 1496 29765 1501 29829
rect 977 29749 1501 29765
rect 977 29685 982 29749
rect 1046 29685 1072 29749
rect 1136 29685 1162 29749
rect 1226 29685 1252 29749
rect 1316 29685 1342 29749
rect 1406 29685 1432 29749
rect 1496 29685 1501 29749
rect 977 29669 1501 29685
rect 977 29605 982 29669
rect 1046 29605 1072 29669
rect 1136 29605 1162 29669
rect 1226 29605 1252 29669
rect 1316 29605 1342 29669
rect 1406 29605 1432 29669
rect 1496 29605 1501 29669
rect 977 29589 1501 29605
rect 977 29525 982 29589
rect 1046 29525 1072 29589
rect 1136 29525 1162 29589
rect 1226 29525 1252 29589
rect 1316 29525 1342 29589
rect 1406 29525 1432 29589
rect 1496 29525 1501 29589
rect 977 29509 1501 29525
rect 977 29445 982 29509
rect 1046 29445 1072 29509
rect 1136 29445 1162 29509
rect 1226 29445 1252 29509
rect 1316 29445 1342 29509
rect 1406 29445 1432 29509
rect 1496 29445 1501 29509
rect 977 29429 1501 29445
rect 977 29365 982 29429
rect 1046 29365 1072 29429
rect 1136 29365 1162 29429
rect 1226 29365 1252 29429
rect 1316 29365 1342 29429
rect 1406 29365 1432 29429
rect 1496 29365 1501 29429
rect 977 29349 1501 29365
rect 977 29285 982 29349
rect 1046 29285 1072 29349
rect 1136 29285 1162 29349
rect 1226 29285 1252 29349
rect 1316 29285 1342 29349
rect 1406 29285 1432 29349
rect 1496 29285 1501 29349
rect 977 29269 1501 29285
rect 977 29205 982 29269
rect 1046 29205 1072 29269
rect 1136 29205 1162 29269
rect 1226 29205 1252 29269
rect 1316 29205 1342 29269
rect 1406 29205 1432 29269
rect 1496 29205 1501 29269
rect 977 29189 1501 29205
rect 977 29125 982 29189
rect 1046 29125 1072 29189
rect 1136 29125 1162 29189
rect 1226 29125 1252 29189
rect 1316 29125 1342 29189
rect 1406 29125 1432 29189
rect 1496 29125 1501 29189
rect 977 29109 1501 29125
rect 977 29045 982 29109
rect 1046 29045 1072 29109
rect 1136 29045 1162 29109
rect 1226 29045 1252 29109
rect 1316 29045 1342 29109
rect 1406 29045 1432 29109
rect 1496 29045 1501 29109
rect 977 29029 1501 29045
rect 977 28965 982 29029
rect 1046 28965 1072 29029
rect 1136 28965 1162 29029
rect 1226 28965 1252 29029
rect 1316 28965 1342 29029
rect 1406 28965 1432 29029
rect 1496 28965 1501 29029
rect 977 28949 1501 28965
rect 977 28885 982 28949
rect 1046 28885 1072 28949
rect 1136 28885 1162 28949
rect 1226 28885 1252 28949
rect 1316 28885 1342 28949
rect 1406 28885 1432 28949
rect 1496 28885 1501 28949
rect 977 28869 1501 28885
rect 977 28805 982 28869
rect 1046 28805 1072 28869
rect 1136 28805 1162 28869
rect 1226 28805 1252 28869
rect 1316 28805 1342 28869
rect 1406 28805 1432 28869
rect 1496 28805 1501 28869
rect 977 28789 1501 28805
rect 977 28725 982 28789
rect 1046 28725 1072 28789
rect 1136 28725 1162 28789
rect 1226 28725 1252 28789
rect 1316 28725 1342 28789
rect 1406 28725 1432 28789
rect 1496 28725 1501 28789
rect 977 28709 1501 28725
rect 977 28645 982 28709
rect 1046 28645 1072 28709
rect 1136 28645 1162 28709
rect 1226 28645 1252 28709
rect 1316 28645 1342 28709
rect 1406 28645 1432 28709
rect 1496 28645 1501 28709
rect 977 28629 1501 28645
rect 977 28565 982 28629
rect 1046 28565 1072 28629
rect 1136 28565 1162 28629
rect 1226 28565 1252 28629
rect 1316 28565 1342 28629
rect 1406 28565 1432 28629
rect 1496 28565 1501 28629
rect 977 28549 1501 28565
rect 977 28485 982 28549
rect 1046 28485 1072 28549
rect 1136 28485 1162 28549
rect 1226 28485 1252 28549
rect 1316 28485 1342 28549
rect 1406 28485 1432 28549
rect 1496 28485 1501 28549
rect 977 28469 1501 28485
rect 977 28405 982 28469
rect 1046 28405 1072 28469
rect 1136 28405 1162 28469
rect 1226 28405 1252 28469
rect 1316 28405 1342 28469
rect 1406 28405 1432 28469
rect 1496 28405 1501 28469
rect 977 28389 1501 28405
rect 977 28325 982 28389
rect 1046 28325 1072 28389
rect 1136 28325 1162 28389
rect 1226 28325 1252 28389
rect 1316 28325 1342 28389
rect 1406 28325 1432 28389
rect 1496 28325 1501 28389
rect 977 28309 1501 28325
rect 977 28245 982 28309
rect 1046 28245 1072 28309
rect 1136 28245 1162 28309
rect 1226 28245 1252 28309
rect 1316 28245 1342 28309
rect 1406 28245 1432 28309
rect 1496 28245 1501 28309
rect 977 28229 1501 28245
rect 977 28165 982 28229
rect 1046 28165 1072 28229
rect 1136 28165 1162 28229
rect 1226 28165 1252 28229
rect 1316 28165 1342 28229
rect 1406 28165 1432 28229
rect 1496 28165 1501 28229
rect 977 28149 1501 28165
rect 977 28085 982 28149
rect 1046 28085 1072 28149
rect 1136 28085 1162 28149
rect 1226 28085 1252 28149
rect 1316 28085 1342 28149
rect 1406 28085 1432 28149
rect 1496 28085 1501 28149
rect 977 28069 1501 28085
rect 977 28005 982 28069
rect 1046 28005 1072 28069
rect 1136 28005 1162 28069
rect 1226 28005 1252 28069
rect 1316 28005 1342 28069
rect 1406 28005 1432 28069
rect 1496 28005 1501 28069
rect 977 27989 1501 28005
rect 977 27925 982 27989
rect 1046 27925 1072 27989
rect 1136 27925 1162 27989
rect 1226 27925 1252 27989
rect 1316 27925 1342 27989
rect 1406 27925 1432 27989
rect 1496 27925 1501 27989
rect 977 27909 1501 27925
rect 977 27845 982 27909
rect 1046 27845 1072 27909
rect 1136 27845 1162 27909
rect 1226 27845 1252 27909
rect 1316 27845 1342 27909
rect 1406 27845 1432 27909
rect 1496 27845 1501 27909
rect 977 27829 1501 27845
rect 977 27765 982 27829
rect 1046 27765 1072 27829
rect 1136 27765 1162 27829
rect 1226 27765 1252 27829
rect 1316 27765 1342 27829
rect 1406 27765 1432 27829
rect 1496 27765 1501 27829
rect 977 27749 1501 27765
rect 977 27685 982 27749
rect 1046 27685 1072 27749
rect 1136 27685 1162 27749
rect 1226 27685 1252 27749
rect 1316 27685 1342 27749
rect 1406 27685 1432 27749
rect 1496 27685 1501 27749
rect 977 27669 1501 27685
rect 977 27605 982 27669
rect 1046 27605 1072 27669
rect 1136 27605 1162 27669
rect 1226 27605 1252 27669
rect 1316 27605 1342 27669
rect 1406 27605 1432 27669
rect 1496 27605 1501 27669
rect 977 27589 1501 27605
rect 977 27525 982 27589
rect 1046 27525 1072 27589
rect 1136 27525 1162 27589
rect 1226 27525 1252 27589
rect 1316 27525 1342 27589
rect 1406 27525 1432 27589
rect 1496 27525 1501 27589
rect 977 27509 1501 27525
rect 977 27445 982 27509
rect 1046 27445 1072 27509
rect 1136 27445 1162 27509
rect 1226 27445 1252 27509
rect 1316 27445 1342 27509
rect 977 27429 1384 27445
rect 977 27365 982 27429
rect 1046 27365 1072 27429
rect 1136 27365 1162 27429
rect 1226 27365 1252 27429
rect 1316 27365 1342 27429
rect 977 27349 1384 27365
rect 977 27285 982 27349
rect 1046 27285 1072 27349
rect 1136 27285 1162 27349
rect 1226 27285 1252 27349
rect 1316 27285 1342 27349
rect 977 27269 1384 27285
rect 977 27205 982 27269
rect 1046 27205 1072 27269
rect 1136 27205 1162 27269
rect 1226 27205 1252 27269
rect 1316 27205 1342 27269
rect 977 27189 1384 27205
rect 977 27125 982 27189
rect 1046 27125 1072 27189
rect 1136 27125 1162 27189
rect 1226 27125 1252 27189
rect 1316 27125 1342 27189
rect 977 27109 1384 27125
rect 977 27045 982 27109
rect 1046 27045 1072 27109
rect 1136 27045 1162 27109
rect 1226 27045 1252 27109
rect 1316 27045 1342 27109
rect 977 27029 1384 27045
rect 977 26965 982 27029
rect 1046 26965 1072 27029
rect 1136 26965 1162 27029
rect 1226 26965 1252 27029
rect 1316 26965 1342 27029
rect 977 26949 1384 26965
rect 977 26885 982 26949
rect 1046 26885 1072 26949
rect 1136 26885 1162 26949
rect 1226 26885 1252 26949
rect 1316 26885 1342 26949
rect 977 26869 1384 26885
rect 977 26805 982 26869
rect 1046 26805 1072 26869
rect 1136 26805 1162 26869
rect 1226 26805 1252 26869
rect 1316 26805 1342 26869
rect 977 26789 1384 26805
rect 977 26725 982 26789
rect 1046 26725 1072 26789
rect 1136 26725 1162 26789
rect 1226 26725 1252 26789
rect 1316 26725 1342 26789
rect 977 26709 1384 26725
rect 977 26645 982 26709
rect 1046 26645 1072 26709
rect 1136 26645 1162 26709
rect 1226 26645 1252 26709
rect 1316 26645 1342 26709
rect 1406 26645 1432 27509
rect 1496 26645 1501 27509
rect 977 26629 1501 26645
rect 977 26565 982 26629
rect 1046 26565 1072 26629
rect 1136 26565 1162 26629
rect 1226 26565 1252 26629
rect 1316 26565 1342 26629
rect 1406 26565 1432 26629
rect 1496 26565 1501 26629
rect 977 26549 1501 26565
rect 977 26485 982 26549
rect 1046 26485 1072 26549
rect 1136 26485 1162 26549
rect 1226 26485 1252 26549
rect 1316 26485 1342 26549
rect 1406 26485 1432 26549
rect 1496 26485 1501 26549
rect 977 26469 1501 26485
rect 977 26405 982 26469
rect 1046 26405 1072 26469
rect 1136 26405 1162 26469
rect 1226 26405 1252 26469
rect 1316 26405 1342 26469
rect 1406 26405 1432 26469
rect 1496 26405 1501 26469
rect 977 26389 1501 26405
rect 977 26325 982 26389
rect 1046 26325 1072 26389
rect 1136 26325 1162 26389
rect 1226 26325 1252 26389
rect 1316 26325 1342 26389
rect 1406 26325 1432 26389
rect 1496 26325 1501 26389
rect 977 26309 1501 26325
rect 977 26245 982 26309
rect 1046 26245 1072 26309
rect 1136 26245 1162 26309
rect 1226 26245 1252 26309
rect 1316 26245 1342 26309
rect 1406 26245 1432 26309
rect 1496 26245 1501 26309
rect 977 26229 1501 26245
rect 977 26165 982 26229
rect 1046 26165 1072 26229
rect 1136 26165 1162 26229
rect 1226 26165 1252 26229
rect 1316 26165 1342 26229
rect 1406 26165 1432 26229
rect 1496 26165 1501 26229
rect 977 26149 1501 26165
rect 977 26085 982 26149
rect 1046 26085 1072 26149
rect 1136 26085 1162 26149
rect 1226 26085 1252 26149
rect 1316 26085 1342 26149
rect 1406 26085 1432 26149
rect 1496 26085 1501 26149
rect 977 26069 1501 26085
rect 977 26005 982 26069
rect 1046 26005 1072 26069
rect 1136 26005 1162 26069
rect 1226 26005 1252 26069
rect 1316 26005 1342 26069
rect 1406 26005 1432 26069
rect 1496 26005 1501 26069
rect 977 25989 1501 26005
rect 977 25925 982 25989
rect 1046 25925 1072 25989
rect 1136 25925 1162 25989
rect 1226 25925 1252 25989
rect 1316 25925 1342 25989
rect 1406 25925 1432 25989
rect 1496 25925 1501 25989
rect 977 25909 1501 25925
rect 977 25845 982 25909
rect 1046 25845 1072 25909
rect 1136 25845 1162 25909
rect 1226 25845 1252 25909
rect 1316 25845 1342 25909
rect 1406 25845 1432 25909
rect 1496 25845 1501 25909
rect 977 25829 1501 25845
rect 977 25765 982 25829
rect 1046 25765 1072 25829
rect 1136 25765 1162 25829
rect 1226 25765 1252 25829
rect 1316 25765 1342 25829
rect 1406 25765 1432 25829
rect 1496 25765 1501 25829
rect 977 25749 1501 25765
rect 977 25685 982 25749
rect 1046 25685 1072 25749
rect 1136 25685 1162 25749
rect 1226 25685 1252 25749
rect 1316 25685 1342 25749
rect 1406 25685 1432 25749
rect 1496 25685 1501 25749
rect 977 25669 1501 25685
rect 977 25605 982 25669
rect 1046 25605 1072 25669
rect 1136 25605 1162 25669
rect 1226 25605 1252 25669
rect 1316 25605 1342 25669
rect 1406 25605 1432 25669
rect 1496 25605 1501 25669
rect 977 25589 1501 25605
rect 977 25525 982 25589
rect 1046 25525 1072 25589
rect 1136 25525 1162 25589
rect 1226 25525 1252 25589
rect 1316 25525 1342 25589
rect 1406 25525 1432 25589
rect 1496 25525 1501 25589
rect 977 25509 1501 25525
rect 977 25445 982 25509
rect 1046 25445 1072 25509
rect 1136 25445 1162 25509
rect 1226 25445 1252 25509
rect 1316 25445 1342 25509
rect 1406 25445 1432 25509
rect 1496 25445 1501 25509
rect 977 25429 1501 25445
rect 977 25365 982 25429
rect 1046 25365 1072 25429
rect 1136 25365 1162 25429
rect 1226 25365 1252 25429
rect 1316 25365 1342 25429
rect 1406 25365 1432 25429
rect 1496 25365 1501 25429
rect 977 25349 1501 25365
rect 977 25285 982 25349
rect 1046 25285 1072 25349
rect 1136 25285 1162 25349
rect 1226 25285 1252 25349
rect 1316 25285 1342 25349
rect 1406 25285 1432 25349
rect 1496 25285 1501 25349
rect 977 25269 1501 25285
rect 977 25205 982 25269
rect 1046 25205 1072 25269
rect 1136 25205 1162 25269
rect 1226 25205 1252 25269
rect 1316 25205 1342 25269
rect 1406 25205 1432 25269
rect 1496 25205 1501 25269
rect 977 25189 1501 25205
rect 977 25125 982 25189
rect 1046 25125 1072 25189
rect 1136 25125 1162 25189
rect 1226 25125 1252 25189
rect 1316 25125 1342 25189
rect 1406 25125 1432 25189
rect 1496 25125 1501 25189
rect 977 25109 1501 25125
rect 977 25045 982 25109
rect 1046 25045 1072 25109
rect 1136 25045 1162 25109
rect 1226 25045 1252 25109
rect 1316 25045 1342 25109
rect 1406 25045 1432 25109
rect 1496 25045 1501 25109
rect 977 25029 1501 25045
rect 977 24965 982 25029
rect 1046 24965 1072 25029
rect 1136 24965 1162 25029
rect 1226 24965 1252 25029
rect 1316 24965 1342 25029
rect 1406 24965 1432 25029
rect 1496 24965 1501 25029
rect 977 24949 1501 24965
rect 977 24885 982 24949
rect 1046 24885 1072 24949
rect 1136 24885 1162 24949
rect 1226 24885 1252 24949
rect 1316 24885 1342 24949
rect 1406 24885 1432 24949
rect 1496 24885 1501 24949
rect 977 24869 1501 24885
rect 977 24805 982 24869
rect 1046 24805 1072 24869
rect 1136 24805 1162 24869
rect 1226 24805 1252 24869
rect 1316 24805 1342 24869
rect 1406 24805 1432 24869
rect 1496 24805 1501 24869
rect 977 24789 1501 24805
rect 977 24725 982 24789
rect 1046 24725 1072 24789
rect 1136 24725 1162 24789
rect 1226 24725 1252 24789
rect 1316 24725 1342 24789
rect 1406 24725 1432 24789
rect 1496 24725 1501 24789
rect 977 24709 1501 24725
rect 977 24645 982 24709
rect 1046 24645 1072 24709
rect 1136 24645 1162 24709
rect 1226 24645 1252 24709
rect 1316 24645 1342 24709
rect 1406 24645 1432 24709
rect 1496 24645 1501 24709
rect 977 24629 1501 24645
rect 977 24565 982 24629
rect 1046 24565 1072 24629
rect 1136 24565 1162 24629
rect 1226 24565 1252 24629
rect 1316 24565 1342 24629
rect 1406 24565 1432 24629
rect 1496 24565 1501 24629
rect 977 24549 1501 24565
rect 977 24485 982 24549
rect 1046 24485 1072 24549
rect 1136 24485 1162 24549
rect 1226 24485 1252 24549
rect 1316 24485 1342 24549
rect 1406 24485 1432 24549
rect 1496 24485 1501 24549
rect 977 24469 1501 24485
rect 977 24405 982 24469
rect 1046 24405 1072 24469
rect 1136 24405 1162 24469
rect 1226 24405 1252 24469
rect 1316 24405 1342 24469
rect 1406 24405 1432 24469
rect 1496 24405 1501 24469
rect 977 24389 1501 24405
rect 977 24325 982 24389
rect 1046 24325 1072 24389
rect 1136 24325 1162 24389
rect 1226 24325 1252 24389
rect 1316 24325 1342 24389
rect 1406 24325 1432 24389
rect 1496 24325 1501 24389
rect 977 24309 1501 24325
rect 977 24245 982 24309
rect 1046 24245 1072 24309
rect 1136 24245 1162 24309
rect 1226 24245 1252 24309
rect 1316 24245 1342 24309
rect 1406 24245 1432 24309
rect 1496 24245 1501 24309
rect 977 24229 1501 24245
rect 977 24165 982 24229
rect 1046 24165 1072 24229
rect 1136 24165 1162 24229
rect 1226 24165 1252 24229
rect 1316 24165 1342 24229
rect 1406 24165 1432 24229
rect 1496 24165 1501 24229
rect 977 24149 1501 24165
rect 977 24085 982 24149
rect 1046 24085 1072 24149
rect 1136 24085 1162 24149
rect 1226 24085 1252 24149
rect 1316 24085 1342 24149
rect 1406 24085 1432 24149
rect 1496 24085 1501 24149
rect 977 24069 1501 24085
rect 977 24005 982 24069
rect 1046 24005 1072 24069
rect 1136 24005 1162 24069
rect 1226 24005 1252 24069
rect 1316 24005 1342 24069
rect 1406 24005 1432 24069
rect 1496 24005 1501 24069
rect 977 23989 1501 24005
rect 977 23925 982 23989
rect 1046 23925 1072 23989
rect 1136 23925 1162 23989
rect 1226 23925 1252 23989
rect 1316 23925 1342 23989
rect 1406 23925 1432 23989
rect 1496 23925 1501 23989
rect 977 23909 1501 23925
rect 977 23845 982 23909
rect 1046 23845 1072 23909
rect 1136 23845 1162 23909
rect 1226 23845 1252 23909
rect 1316 23845 1342 23909
rect 1406 23845 1432 23909
rect 1496 23845 1501 23909
rect 977 23829 1501 23845
rect 977 23765 982 23829
rect 1046 23765 1072 23829
rect 1136 23765 1162 23829
rect 1226 23765 1252 23829
rect 1316 23765 1342 23829
rect 1406 23765 1432 23829
rect 1496 23765 1501 23829
rect 977 23749 1501 23765
rect 977 23685 982 23749
rect 1046 23685 1072 23749
rect 1136 23685 1162 23749
rect 1226 23685 1252 23749
rect 1316 23685 1342 23749
rect 1406 23685 1432 23749
rect 1496 23685 1501 23749
rect 977 23669 1501 23685
rect 977 23605 982 23669
rect 1046 23605 1072 23669
rect 1136 23605 1162 23669
rect 1226 23605 1252 23669
rect 1316 23605 1342 23669
rect 1406 23605 1432 23669
rect 1496 23605 1501 23669
rect 977 23589 1501 23605
rect 977 23525 982 23589
rect 1046 23525 1072 23589
rect 1136 23525 1162 23589
rect 1226 23525 1252 23589
rect 1316 23525 1342 23589
rect 1406 23525 1432 23589
rect 1496 23525 1501 23589
rect 977 23509 1501 23525
rect 977 23445 982 23509
rect 1046 23445 1072 23509
rect 1136 23445 1162 23509
rect 1226 23445 1252 23509
rect 1316 23445 1342 23509
rect 1406 23445 1432 23509
rect 1496 23445 1501 23509
rect 977 23429 1501 23445
rect 977 23365 982 23429
rect 1046 23365 1072 23429
rect 1136 23365 1162 23429
rect 1226 23365 1252 23429
rect 1316 23365 1342 23429
rect 1406 23365 1432 23429
rect 1496 23365 1501 23429
rect 977 23349 1501 23365
rect 977 23285 982 23349
rect 1046 23285 1072 23349
rect 1136 23285 1162 23349
rect 1226 23285 1252 23349
rect 1316 23285 1342 23349
rect 1406 23285 1432 23349
rect 1496 23285 1501 23349
rect 977 23268 1501 23285
rect 977 23204 982 23268
rect 1046 23204 1072 23268
rect 1136 23204 1162 23268
rect 1226 23204 1252 23268
rect 1316 23204 1342 23268
rect 1406 23204 1432 23268
rect 1496 23204 1501 23268
rect 977 23187 1501 23204
rect 977 23123 982 23187
rect 1046 23123 1072 23187
rect 1136 23123 1162 23187
rect 1226 23123 1252 23187
rect 1316 23123 1342 23187
rect 1406 23123 1432 23187
rect 1496 23123 1501 23187
rect 977 23106 1501 23123
rect 977 23042 982 23106
rect 1046 23042 1072 23106
rect 1136 23042 1162 23106
rect 1226 23042 1252 23106
rect 1316 23042 1342 23106
rect 1406 23042 1432 23106
rect 1496 23042 1501 23106
rect 977 23025 1501 23042
rect 977 22961 982 23025
rect 1046 22961 1072 23025
rect 1136 22961 1162 23025
rect 1226 22961 1252 23025
rect 1316 22961 1342 23025
rect 1406 22961 1432 23025
rect 1496 22961 1501 23025
rect 977 22944 1501 22961
rect 977 22880 982 22944
rect 1046 22880 1072 22944
rect 1136 22880 1162 22944
rect 1226 22880 1252 22944
rect 1316 22880 1342 22944
rect 1406 22880 1432 22944
rect 1496 22880 1501 22944
rect 977 22863 1501 22880
rect 977 22799 982 22863
rect 1046 22799 1072 22863
rect 1136 22799 1162 22863
rect 1226 22799 1252 22863
rect 1316 22799 1342 22863
rect 1406 22799 1432 22863
rect 1496 22799 1501 22863
rect 977 22782 1501 22799
rect 977 22718 982 22782
rect 1046 22718 1072 22782
rect 1136 22718 1162 22782
rect 1226 22718 1252 22782
rect 1316 22718 1342 22782
rect 1406 22718 1432 22782
rect 1496 22718 1501 22782
rect 977 22701 1501 22718
rect 977 22637 982 22701
rect 1046 22637 1072 22701
rect 1136 22637 1162 22701
rect 1226 22637 1252 22701
rect 1316 22637 1342 22701
rect 1406 22637 1432 22701
rect 1496 22637 1501 22701
rect 977 22620 1501 22637
rect 977 22556 982 22620
rect 1046 22556 1072 22620
rect 1136 22556 1162 22620
rect 1226 22556 1252 22620
rect 1316 22556 1342 22620
rect 1406 22556 1432 22620
rect 1496 22556 1501 22620
rect 977 22539 1501 22556
rect 977 22475 982 22539
rect 1046 22475 1072 22539
rect 1136 22475 1162 22539
rect 1226 22475 1252 22539
rect 1316 22475 1342 22539
rect 1406 22475 1432 22539
rect 1496 22475 1501 22539
rect 977 22458 1501 22475
rect 977 22394 982 22458
rect 1046 22394 1072 22458
rect 1136 22394 1162 22458
rect 1226 22394 1252 22458
rect 1316 22394 1342 22458
rect 1406 22394 1432 22458
rect 1496 22394 1501 22458
rect 977 22377 1501 22394
rect 977 22313 982 22377
rect 1046 22313 1072 22377
rect 1136 22313 1162 22377
rect 1226 22313 1252 22377
rect 1316 22313 1342 22377
rect 1406 22313 1432 22377
rect 1496 22313 1501 22377
rect 977 22296 1501 22313
rect 977 22232 982 22296
rect 1046 22232 1072 22296
rect 1136 22232 1162 22296
rect 1226 22232 1252 22296
rect 1316 22232 1342 22296
rect 1406 22232 1432 22296
rect 1496 22232 1501 22296
rect 977 22215 1501 22232
rect 977 22151 982 22215
rect 1046 22151 1072 22215
rect 1136 22151 1162 22215
rect 1226 22151 1252 22215
rect 1316 22151 1342 22215
rect 1406 22151 1432 22215
rect 1496 22151 1501 22215
rect 977 22134 1501 22151
rect 977 22070 982 22134
rect 1046 22070 1072 22134
rect 1136 22070 1162 22134
rect 1226 22070 1252 22134
rect 1316 22070 1342 22134
rect 1406 22070 1432 22134
rect 1496 22070 1501 22134
rect 977 22053 1501 22070
rect 977 21989 982 22053
rect 1046 21989 1072 22053
rect 1136 21989 1162 22053
rect 1226 21989 1252 22053
rect 1316 21989 1342 22053
rect 1406 21989 1432 22053
rect 1496 21989 1501 22053
rect 977 21972 1501 21989
rect 977 21908 982 21972
rect 1046 21908 1072 21972
rect 1136 21908 1162 21972
rect 1226 21908 1252 21972
rect 1316 21908 1342 21972
rect 1406 21908 1432 21972
rect 1496 21908 1501 21972
rect 977 21891 1501 21908
rect 977 21827 982 21891
rect 1046 21827 1072 21891
rect 1136 21827 1162 21891
rect 1226 21827 1252 21891
rect 1316 21827 1342 21891
rect 1406 21827 1432 21891
rect 1496 21827 1501 21891
rect 977 21810 1501 21827
rect 977 21746 982 21810
rect 1046 21746 1072 21810
rect 1136 21746 1162 21810
rect 1226 21746 1252 21810
rect 1316 21746 1342 21810
rect 1406 21746 1432 21810
rect 1496 21746 1501 21810
rect 977 21729 1501 21746
rect 977 21665 982 21729
rect 1046 21665 1072 21729
rect 1136 21665 1162 21729
rect 1226 21665 1252 21729
rect 1316 21665 1342 21729
rect 1406 21665 1432 21729
rect 1496 21665 1501 21729
rect 977 21648 1501 21665
rect 977 21584 982 21648
rect 1046 21584 1072 21648
rect 1136 21584 1162 21648
rect 1226 21584 1252 21648
rect 1316 21584 1342 21648
rect 1406 21584 1432 21648
rect 1496 21584 1501 21648
rect 977 21567 1501 21584
rect 977 21503 982 21567
rect 1046 21503 1072 21567
rect 1136 21503 1162 21567
rect 1226 21503 1252 21567
rect 1316 21503 1342 21567
rect 1406 21503 1432 21567
rect 1496 21503 1501 21567
rect 977 21486 1501 21503
rect 977 21422 982 21486
rect 1046 21422 1072 21486
rect 1136 21422 1162 21486
rect 1226 21422 1252 21486
rect 1316 21422 1342 21486
rect 1406 21422 1432 21486
rect 1496 21422 1501 21486
rect 977 21405 1501 21422
rect 977 21341 982 21405
rect 1046 21341 1072 21405
rect 1136 21341 1162 21405
rect 1226 21341 1252 21405
rect 1316 21341 1342 21405
rect 1406 21341 1432 21405
rect 1496 21341 1501 21405
rect 977 21324 1501 21341
rect 977 21260 982 21324
rect 1046 21260 1072 21324
rect 1136 21260 1162 21324
rect 1226 21260 1252 21324
rect 1316 21260 1342 21324
rect 1406 21260 1432 21324
rect 1496 21260 1501 21324
rect 977 21243 1501 21260
rect 977 21179 982 21243
rect 1046 21179 1072 21243
rect 1136 21179 1162 21243
rect 1226 21179 1252 21243
rect 1316 21179 1342 21243
rect 1406 21179 1432 21243
rect 1496 21179 1501 21243
rect 977 21162 1501 21179
rect 977 21098 982 21162
rect 1046 21098 1072 21162
rect 1136 21098 1162 21162
rect 1226 21098 1252 21162
rect 1316 21098 1342 21162
rect 1406 21098 1432 21162
rect 1496 21098 1501 21162
rect 977 21081 1501 21098
rect 977 21017 982 21081
rect 1046 21017 1072 21081
rect 1136 21017 1162 21081
rect 1226 21017 1252 21081
rect 1316 21017 1342 21081
rect 1406 21017 1432 21081
rect 1496 21017 1501 21081
rect 977 21000 1501 21017
rect 977 20936 982 21000
rect 1046 20936 1072 21000
rect 1136 20936 1162 21000
rect 1226 20936 1252 21000
rect 1316 20936 1342 21000
rect 1406 20936 1432 21000
rect 1496 20972 1501 21000
rect 13515 33109 14039 33110
rect 13515 33045 13520 33109
rect 13584 33045 13610 33109
rect 13674 33045 13700 33109
rect 13764 33045 13790 33109
rect 13854 33045 13880 33109
rect 13944 33045 13970 33109
rect 14034 33045 14039 33109
rect 13515 33029 14039 33045
rect 13515 32965 13520 33029
rect 13584 32965 13610 33029
rect 13674 32965 13700 33029
rect 13764 32965 13790 33029
rect 13854 32965 13880 33029
rect 13944 32965 13970 33029
rect 14034 32965 14039 33029
rect 13515 32949 14039 32965
rect 13515 32885 13520 32949
rect 13584 32885 13610 32949
rect 13674 32885 13700 32949
rect 13764 32885 13790 32949
rect 13854 32885 13880 32949
rect 13944 32885 13970 32949
rect 14034 32885 14039 32949
rect 13515 32869 14039 32885
rect 13515 32805 13520 32869
rect 13584 32805 13610 32869
rect 13674 32805 13700 32869
rect 13764 32805 13790 32869
rect 13854 32805 13880 32869
rect 13944 32805 13970 32869
rect 14034 32805 14039 32869
rect 13515 32789 14039 32805
rect 13515 32725 13520 32789
rect 13584 32725 13610 32789
rect 13674 32725 13700 32789
rect 13764 32725 13790 32789
rect 13854 32725 13880 32789
rect 13944 32725 13970 32789
rect 14034 32725 14039 32789
rect 13515 32709 14039 32725
rect 13515 32645 13520 32709
rect 13584 32645 13610 32709
rect 13674 32645 13700 32709
rect 13764 32645 13790 32709
rect 13854 32645 13880 32709
rect 13944 32645 13970 32709
rect 14034 32645 14039 32709
rect 13515 32629 14039 32645
rect 13515 32565 13520 32629
rect 13584 32565 13610 32629
rect 13674 32565 13700 32629
rect 13764 32565 13790 32629
rect 13854 32565 13880 32629
rect 13944 32565 13970 32629
rect 14034 32565 14039 32629
rect 13515 32549 14039 32565
rect 13515 32485 13520 32549
rect 13584 32485 13610 32549
rect 13674 32485 13700 32549
rect 13764 32485 13790 32549
rect 13854 32485 13880 32549
rect 13944 32485 13970 32549
rect 14034 32485 14039 32549
rect 13515 32469 14039 32485
rect 13515 32405 13520 32469
rect 13584 32405 13610 32469
rect 13674 32405 13700 32469
rect 13764 32405 13790 32469
rect 13854 32405 13880 32469
rect 13944 32405 13970 32469
rect 14034 32405 14039 32469
rect 13515 32389 14039 32405
rect 13515 32325 13520 32389
rect 13584 32325 13610 32389
rect 13674 32325 13700 32389
rect 13764 32325 13790 32389
rect 13854 32325 13880 32389
rect 13944 32325 13970 32389
rect 14034 32325 14039 32389
rect 13515 32309 14039 32325
rect 13515 32245 13520 32309
rect 13584 32245 13610 32309
rect 13674 32245 13700 32309
rect 13764 32245 13790 32309
rect 13854 32245 13880 32309
rect 13944 32245 13970 32309
rect 14034 32245 14039 32309
rect 13515 32229 14039 32245
rect 13515 32165 13520 32229
rect 13584 32165 13610 32229
rect 13674 32165 13700 32229
rect 13764 32165 13790 32229
rect 13854 32165 13880 32229
rect 13944 32165 13970 32229
rect 14034 32165 14039 32229
rect 13515 32149 14039 32165
rect 13515 32085 13520 32149
rect 13584 32085 13610 32149
rect 13674 32085 13700 32149
rect 13764 32085 13790 32149
rect 13854 32085 13880 32149
rect 13944 32085 13970 32149
rect 14034 32085 14039 32149
rect 13515 32069 14039 32085
rect 13515 32005 13520 32069
rect 13584 32005 13610 32069
rect 13674 32005 13700 32069
rect 13764 32005 13790 32069
rect 13854 32005 13880 32069
rect 13944 32005 13970 32069
rect 14034 32005 14039 32069
rect 13515 31989 14039 32005
rect 13515 31925 13520 31989
rect 13584 31925 13610 31989
rect 13674 31925 13700 31989
rect 13764 31925 13790 31989
rect 13854 31925 13880 31989
rect 13944 31925 13970 31989
rect 14034 31925 14039 31989
rect 13515 31909 14039 31925
rect 13515 31845 13520 31909
rect 13584 31845 13610 31909
rect 13674 31845 13700 31909
rect 13764 31845 13790 31909
rect 13854 31845 13880 31909
rect 13944 31845 13970 31909
rect 14034 31845 14039 31909
rect 13515 31829 14039 31845
rect 13515 31765 13520 31829
rect 13584 31765 13610 31829
rect 13674 31765 13700 31829
rect 13764 31765 13790 31829
rect 13854 31765 13880 31829
rect 13944 31765 13970 31829
rect 14034 31765 14039 31829
rect 13515 31749 14039 31765
rect 13515 31685 13520 31749
rect 13584 31685 13610 31749
rect 13674 31685 13700 31749
rect 13764 31685 13790 31749
rect 13854 31685 13880 31749
rect 13944 31685 13970 31749
rect 14034 31685 14039 31749
rect 13515 31669 14039 31685
rect 13515 31605 13520 31669
rect 13584 31605 13610 31669
rect 13674 31605 13700 31669
rect 13764 31605 13790 31669
rect 13854 31605 13880 31669
rect 13944 31605 13970 31669
rect 14034 31605 14039 31669
rect 13515 31589 14039 31605
rect 13515 31525 13520 31589
rect 13584 31525 13610 31589
rect 13674 31525 13700 31589
rect 13764 31525 13790 31589
rect 13854 31525 13880 31589
rect 13944 31525 13970 31589
rect 14034 31525 14039 31589
rect 13515 31509 14039 31525
rect 13515 31445 13520 31509
rect 13584 31445 13610 31509
rect 13674 31445 13700 31509
rect 13764 31445 13790 31509
rect 13854 31445 13880 31509
rect 13944 31445 13970 31509
rect 14034 31445 14039 31509
rect 13515 31429 14039 31445
rect 13515 31365 13520 31429
rect 13584 31365 13610 31429
rect 13674 31365 13700 31429
rect 13764 31365 13790 31429
rect 13854 31365 13880 31429
rect 13944 31365 13970 31429
rect 14034 31365 14039 31429
rect 13515 31349 14039 31365
rect 13515 31285 13520 31349
rect 13584 31285 13610 31349
rect 13674 31285 13700 31349
rect 13764 31285 13790 31349
rect 13854 31285 13880 31349
rect 13944 31285 13970 31349
rect 14034 31285 14039 31349
rect 13515 31269 14039 31285
rect 13515 31205 13520 31269
rect 13584 31205 13610 31269
rect 13674 31205 13700 31269
rect 13764 31205 13790 31269
rect 13854 31205 13880 31269
rect 13944 31205 13970 31269
rect 14034 31205 14039 31269
rect 13515 31189 14039 31205
rect 13515 31125 13520 31189
rect 13584 31125 13610 31189
rect 13674 31125 13700 31189
rect 13764 31125 13790 31189
rect 13854 31125 13880 31189
rect 13944 31125 13970 31189
rect 14034 31125 14039 31189
rect 13515 31109 14039 31125
rect 13515 31045 13520 31109
rect 13584 31045 13610 31109
rect 13674 31045 13700 31109
rect 13764 31045 13790 31109
rect 13854 31045 13880 31109
rect 13944 31045 13970 31109
rect 14034 31045 14039 31109
rect 13515 31029 14039 31045
rect 13515 30965 13520 31029
rect 13584 30965 13610 31029
rect 13674 30965 13700 31029
rect 13764 30965 13790 31029
rect 13854 30965 13880 31029
rect 13944 30965 13970 31029
rect 14034 30965 14039 31029
rect 13515 30949 14039 30965
rect 13515 30885 13520 30949
rect 13584 30885 13610 30949
rect 13674 30885 13700 30949
rect 13764 30885 13790 30949
rect 13854 30885 13880 30949
rect 13944 30885 13970 30949
rect 14034 30885 14039 30949
rect 13515 30869 14039 30885
rect 13515 30805 13520 30869
rect 13584 30805 13610 30869
rect 13674 30805 13700 30869
rect 13764 30805 13790 30869
rect 13854 30805 13880 30869
rect 13944 30805 13970 30869
rect 14034 30805 14039 30869
rect 13515 30789 14039 30805
rect 13515 30725 13520 30789
rect 13584 30725 13610 30789
rect 13674 30725 13700 30789
rect 13764 30725 13790 30789
rect 13854 30725 13880 30789
rect 13944 30725 13970 30789
rect 14034 30725 14039 30789
rect 13515 30709 14039 30725
rect 13515 30645 13520 30709
rect 13584 30645 13610 30709
rect 13674 30645 13700 30709
rect 13764 30645 13790 30709
rect 13854 30645 13880 30709
rect 13944 30645 13970 30709
rect 14034 30645 14039 30709
rect 13515 30629 14039 30645
rect 13515 30565 13520 30629
rect 13584 30565 13610 30629
rect 13674 30565 13700 30629
rect 13764 30565 13790 30629
rect 13854 30565 13880 30629
rect 13944 30565 13970 30629
rect 14034 30565 14039 30629
rect 13515 30549 14039 30565
rect 13515 30485 13520 30549
rect 13584 30485 13610 30549
rect 13674 30485 13700 30549
rect 13764 30485 13790 30549
rect 13854 30485 13880 30549
rect 13944 30485 13970 30549
rect 14034 30485 14039 30549
rect 13515 30469 14039 30485
rect 13515 30405 13520 30469
rect 13584 30405 13610 30469
rect 13674 30405 13700 30469
rect 13764 30405 13790 30469
rect 13854 30405 13880 30469
rect 13944 30405 13970 30469
rect 14034 30405 14039 30469
rect 13515 30389 14039 30405
rect 13515 30325 13520 30389
rect 13584 30325 13610 30389
rect 13674 30325 13700 30389
rect 13764 30325 13790 30389
rect 13854 30325 13880 30389
rect 13944 30325 13970 30389
rect 14034 30325 14039 30389
rect 13515 30309 14039 30325
rect 13515 30245 13520 30309
rect 13584 30245 13610 30309
rect 13674 30245 13700 30309
rect 13764 30245 13790 30309
rect 13854 30245 13880 30309
rect 13944 30245 13970 30309
rect 14034 30245 14039 30309
rect 13515 30229 14039 30245
rect 13515 30165 13520 30229
rect 13584 30165 13610 30229
rect 13674 30165 13700 30229
rect 13764 30165 13790 30229
rect 13854 30165 13880 30229
rect 13944 30165 13970 30229
rect 14034 30165 14039 30229
rect 13515 30149 14039 30165
rect 13515 30085 13520 30149
rect 13584 30085 13610 30149
rect 13674 30085 13700 30149
rect 13764 30085 13790 30149
rect 13854 30085 13880 30149
rect 13944 30085 13970 30149
rect 14034 30085 14039 30149
rect 13515 30069 14039 30085
rect 13515 30005 13520 30069
rect 13584 30005 13610 30069
rect 13674 30005 13700 30069
rect 13764 30005 13790 30069
rect 13854 30005 13880 30069
rect 13944 30005 13970 30069
rect 14034 30005 14039 30069
rect 13515 29989 14039 30005
rect 13515 29925 13520 29989
rect 13584 29925 13610 29989
rect 13674 29925 13700 29989
rect 13764 29925 13790 29989
rect 13854 29925 13880 29989
rect 13944 29925 13970 29989
rect 14034 29925 14039 29989
rect 13515 29909 14039 29925
rect 13515 29845 13520 29909
rect 13584 29845 13610 29909
rect 13674 29845 13700 29909
rect 13764 29845 13790 29909
rect 13854 29845 13880 29909
rect 13944 29845 13970 29909
rect 14034 29845 14039 29909
rect 13515 29829 14039 29845
rect 13515 29765 13520 29829
rect 13584 29765 13610 29829
rect 13674 29765 13700 29829
rect 13764 29765 13790 29829
rect 13854 29765 13880 29829
rect 13944 29765 13970 29829
rect 14034 29765 14039 29829
rect 13515 29749 14039 29765
rect 13515 29685 13520 29749
rect 13584 29685 13610 29749
rect 13674 29685 13700 29749
rect 13764 29685 13790 29749
rect 13854 29685 13880 29749
rect 13944 29685 13970 29749
rect 14034 29685 14039 29749
rect 13515 29669 14039 29685
rect 13515 29605 13520 29669
rect 13584 29605 13610 29669
rect 13674 29605 13700 29669
rect 13764 29605 13790 29669
rect 13854 29605 13880 29669
rect 13944 29605 13970 29669
rect 14034 29605 14039 29669
rect 13515 29589 14039 29605
rect 13515 29525 13520 29589
rect 13584 29525 13610 29589
rect 13674 29525 13700 29589
rect 13764 29525 13790 29589
rect 13854 29525 13880 29589
rect 13944 29525 13970 29589
rect 14034 29525 14039 29589
rect 13515 29509 14039 29525
rect 13515 29445 13520 29509
rect 13584 29445 13610 29509
rect 13674 29445 13700 29509
rect 13764 29445 13790 29509
rect 13854 29445 13880 29509
rect 13944 29445 13970 29509
rect 14034 29445 14039 29509
rect 13515 29429 14039 29445
rect 13515 29365 13520 29429
rect 13584 29365 13610 29429
rect 13674 29365 13700 29429
rect 13764 29365 13790 29429
rect 13854 29365 13880 29429
rect 13944 29365 13970 29429
rect 14034 29365 14039 29429
rect 13515 29349 14039 29365
rect 13515 29285 13520 29349
rect 13584 29285 13610 29349
rect 13674 29285 13700 29349
rect 13764 29285 13790 29349
rect 13854 29285 13880 29349
rect 13944 29285 13970 29349
rect 14034 29285 14039 29349
rect 13515 29269 14039 29285
rect 13515 29205 13520 29269
rect 13584 29205 13610 29269
rect 13674 29205 13700 29269
rect 13764 29205 13790 29269
rect 13854 29205 13880 29269
rect 13944 29205 13970 29269
rect 14034 29205 14039 29269
rect 13515 29189 14039 29205
rect 13515 29125 13520 29189
rect 13584 29125 13610 29189
rect 13674 29125 13700 29189
rect 13764 29125 13790 29189
rect 13854 29125 13880 29189
rect 13944 29125 13970 29189
rect 14034 29125 14039 29189
rect 13515 29109 14039 29125
rect 13515 29045 13520 29109
rect 13584 29045 13610 29109
rect 13674 29045 13700 29109
rect 13764 29045 13790 29109
rect 13854 29045 13880 29109
rect 13944 29045 13970 29109
rect 14034 29045 14039 29109
rect 13515 29029 14039 29045
rect 13515 28965 13520 29029
rect 13584 28965 13610 29029
rect 13674 28965 13700 29029
rect 13764 28965 13790 29029
rect 13854 28965 13880 29029
rect 13944 28965 13970 29029
rect 14034 28965 14039 29029
rect 13515 28949 14039 28965
rect 13515 28885 13520 28949
rect 13584 28885 13610 28949
rect 13674 28885 13700 28949
rect 13764 28885 13790 28949
rect 13854 28885 13880 28949
rect 13944 28885 13970 28949
rect 14034 28885 14039 28949
rect 13515 28869 14039 28885
rect 13515 28805 13520 28869
rect 13584 28805 13610 28869
rect 13674 28805 13700 28869
rect 13764 28805 13790 28869
rect 13854 28805 13880 28869
rect 13944 28805 13970 28869
rect 14034 28805 14039 28869
rect 13515 28789 14039 28805
rect 13515 28725 13520 28789
rect 13584 28725 13610 28789
rect 13674 28725 13700 28789
rect 13764 28725 13790 28789
rect 13854 28725 13880 28789
rect 13944 28725 13970 28789
rect 14034 28725 14039 28789
rect 13515 28709 14039 28725
rect 13515 28645 13520 28709
rect 13584 28645 13610 28709
rect 13674 28645 13700 28709
rect 13764 28645 13790 28709
rect 13854 28645 13880 28709
rect 13944 28645 13970 28709
rect 14034 28645 14039 28709
rect 13515 28629 14039 28645
rect 13515 28565 13520 28629
rect 13584 28565 13610 28629
rect 13674 28565 13700 28629
rect 13764 28565 13790 28629
rect 13854 28565 13880 28629
rect 13944 28565 13970 28629
rect 14034 28565 14039 28629
rect 13515 28549 14039 28565
rect 13515 28485 13520 28549
rect 13584 28485 13610 28549
rect 13674 28485 13700 28549
rect 13764 28485 13790 28549
rect 13854 28485 13880 28549
rect 13944 28485 13970 28549
rect 14034 28485 14039 28549
rect 13515 28469 14039 28485
rect 13515 28405 13520 28469
rect 13584 28405 13610 28469
rect 13674 28405 13700 28469
rect 13764 28405 13790 28469
rect 13854 28405 13880 28469
rect 13944 28405 13970 28469
rect 14034 28405 14039 28469
rect 13515 28389 14039 28405
rect 13515 28325 13520 28389
rect 13584 28325 13610 28389
rect 13674 28325 13700 28389
rect 13764 28325 13790 28389
rect 13854 28325 13880 28389
rect 13944 28325 13970 28389
rect 14034 28325 14039 28389
rect 13515 28309 14039 28325
rect 13515 28245 13520 28309
rect 13584 28245 13610 28309
rect 13674 28245 13700 28309
rect 13764 28245 13790 28309
rect 13854 28245 13880 28309
rect 13944 28245 13970 28309
rect 14034 28245 14039 28309
rect 13515 28229 14039 28245
rect 13515 28165 13520 28229
rect 13584 28165 13610 28229
rect 13674 28165 13700 28229
rect 13764 28165 13790 28229
rect 13854 28165 13880 28229
rect 13944 28165 13970 28229
rect 14034 28165 14039 28229
rect 13515 28149 14039 28165
rect 13515 28085 13520 28149
rect 13584 28085 13610 28149
rect 13674 28085 13700 28149
rect 13764 28085 13790 28149
rect 13854 28085 13880 28149
rect 13944 28085 13970 28149
rect 14034 28085 14039 28149
rect 13515 28069 14039 28085
rect 13515 28005 13520 28069
rect 13584 28005 13610 28069
rect 13674 28005 13700 28069
rect 13764 28005 13790 28069
rect 13854 28005 13880 28069
rect 13944 28005 13970 28069
rect 14034 28005 14039 28069
rect 13515 27989 14039 28005
rect 13515 27925 13520 27989
rect 13584 27925 13610 27989
rect 13674 27925 13700 27989
rect 13764 27925 13790 27989
rect 13854 27925 13880 27989
rect 13944 27925 13970 27989
rect 14034 27925 14039 27989
rect 13515 27909 14039 27925
rect 13515 27845 13520 27909
rect 13584 27845 13610 27909
rect 13674 27845 13700 27909
rect 13764 27845 13790 27909
rect 13854 27845 13880 27909
rect 13944 27845 13970 27909
rect 14034 27845 14039 27909
rect 13515 27829 14039 27845
rect 13515 27765 13520 27829
rect 13584 27765 13610 27829
rect 13674 27765 13700 27829
rect 13764 27765 13790 27829
rect 13854 27765 13880 27829
rect 13944 27765 13970 27829
rect 14034 27765 14039 27829
rect 13515 27749 14039 27765
rect 13515 27685 13520 27749
rect 13584 27685 13610 27749
rect 13674 27685 13700 27749
rect 13764 27685 13790 27749
rect 13854 27685 13880 27749
rect 13944 27685 13970 27749
rect 14034 27685 14039 27749
rect 13515 27669 14039 27685
rect 13515 27605 13520 27669
rect 13584 27605 13610 27669
rect 13674 27605 13700 27669
rect 13764 27605 13790 27669
rect 13854 27605 13880 27669
rect 13944 27605 13970 27669
rect 14034 27605 14039 27669
rect 13515 27589 14039 27605
rect 13515 27525 13520 27589
rect 13584 27525 13610 27589
rect 13674 27525 13700 27589
rect 13764 27525 13790 27589
rect 13854 27525 13880 27589
rect 13944 27525 13970 27589
rect 14034 27525 14039 27589
rect 13515 27509 14039 27525
rect 13515 27445 13520 27509
rect 13584 27445 13610 27509
rect 13674 27445 13700 27509
rect 13764 27445 13790 27509
rect 13854 27445 13880 27509
rect 13944 27445 13970 27509
rect 14034 27445 14039 27509
rect 13515 27429 14039 27445
rect 13515 27365 13520 27429
rect 13584 27365 13610 27429
rect 13674 27365 13700 27429
rect 13764 27365 13790 27429
rect 13854 27365 13880 27429
rect 13944 27365 13970 27429
rect 14034 27365 14039 27429
rect 13515 27349 14039 27365
rect 13515 27285 13520 27349
rect 13584 27285 13610 27349
rect 13674 27285 13700 27349
rect 13764 27285 13790 27349
rect 13854 27285 13880 27349
rect 13944 27285 13970 27349
rect 14034 27285 14039 27349
rect 13515 27269 14039 27285
rect 13515 27205 13520 27269
rect 13584 27205 13610 27269
rect 13674 27205 13700 27269
rect 13764 27205 13790 27269
rect 13854 27205 13880 27269
rect 13944 27205 13970 27269
rect 14034 27205 14039 27269
rect 13515 27189 14039 27205
rect 13515 27125 13520 27189
rect 13584 27125 13610 27189
rect 13674 27125 13700 27189
rect 13764 27125 13790 27189
rect 13854 27125 13880 27189
rect 13944 27125 13970 27189
rect 14034 27125 14039 27189
rect 13515 27109 14039 27125
rect 13515 27045 13520 27109
rect 13584 27045 13610 27109
rect 13674 27045 13700 27109
rect 13764 27045 13790 27109
rect 13854 27045 13880 27109
rect 13944 27045 13970 27109
rect 14034 27045 14039 27109
rect 13515 27029 14039 27045
rect 13515 26965 13520 27029
rect 13584 26965 13610 27029
rect 13674 26965 13700 27029
rect 13764 26965 13790 27029
rect 13854 26965 13880 27029
rect 13944 26965 13970 27029
rect 14034 26965 14039 27029
rect 13515 26949 14039 26965
rect 13515 26885 13520 26949
rect 13584 26885 13610 26949
rect 13674 26885 13700 26949
rect 13764 26885 13790 26949
rect 13854 26885 13880 26949
rect 13944 26885 13970 26949
rect 14034 26885 14039 26949
rect 13515 26869 14039 26885
rect 13515 26805 13520 26869
rect 13584 26805 13610 26869
rect 13674 26805 13700 26869
rect 13764 26805 13790 26869
rect 13854 26805 13880 26869
rect 13944 26805 13970 26869
rect 14034 26805 14039 26869
rect 13515 26789 14039 26805
rect 13515 26725 13520 26789
rect 13584 26725 13610 26789
rect 13674 26725 13700 26789
rect 13764 26725 13790 26789
rect 13854 26725 13880 26789
rect 13944 26725 13970 26789
rect 14034 26725 14039 26789
rect 13515 26709 14039 26725
rect 13515 26645 13520 26709
rect 13584 26645 13610 26709
rect 13674 26645 13700 26709
rect 13764 26645 13790 26709
rect 13854 26645 13880 26709
rect 13944 26645 13970 26709
rect 14034 26645 14039 26709
rect 13515 26629 14039 26645
rect 13515 26565 13520 26629
rect 13584 26565 13610 26629
rect 13674 26565 13700 26629
rect 13764 26565 13790 26629
rect 13854 26565 13880 26629
rect 13944 26565 13970 26629
rect 14034 26565 14039 26629
rect 13515 26549 14039 26565
rect 13515 26485 13520 26549
rect 13584 26485 13610 26549
rect 13674 26485 13700 26549
rect 13764 26485 13790 26549
rect 13854 26485 13880 26549
rect 13944 26485 13970 26549
rect 14034 26485 14039 26549
rect 13515 26469 14039 26485
rect 13515 26405 13520 26469
rect 13584 26405 13610 26469
rect 13674 26405 13700 26469
rect 13764 26405 13790 26469
rect 13854 26405 13880 26469
rect 13944 26405 13970 26469
rect 14034 26405 14039 26469
rect 13515 26389 14039 26405
rect 13515 26325 13520 26389
rect 13584 26325 13610 26389
rect 13674 26325 13700 26389
rect 13764 26325 13790 26389
rect 13854 26325 13880 26389
rect 13944 26325 13970 26389
rect 14034 26325 14039 26389
rect 13515 26309 14039 26325
rect 13515 26245 13520 26309
rect 13584 26245 13610 26309
rect 13674 26245 13700 26309
rect 13764 26245 13790 26309
rect 13854 26245 13880 26309
rect 13944 26245 13970 26309
rect 14034 26245 14039 26309
rect 13515 26229 14039 26245
rect 13515 26165 13520 26229
rect 13584 26165 13610 26229
rect 13674 26165 13700 26229
rect 13764 26165 13790 26229
rect 13854 26165 13880 26229
rect 13944 26165 13970 26229
rect 14034 26165 14039 26229
rect 13515 26149 14039 26165
rect 13515 26085 13520 26149
rect 13584 26085 13610 26149
rect 13674 26085 13700 26149
rect 13764 26085 13790 26149
rect 13854 26085 13880 26149
rect 13944 26085 13970 26149
rect 14034 26085 14039 26149
rect 13515 26069 14039 26085
rect 13515 26005 13520 26069
rect 13584 26005 13610 26069
rect 13674 26005 13700 26069
rect 13764 26005 13790 26069
rect 13854 26005 13880 26069
rect 13944 26005 13970 26069
rect 14034 26005 14039 26069
rect 13515 25989 14039 26005
rect 13515 25925 13520 25989
rect 13584 25925 13610 25989
rect 13674 25925 13700 25989
rect 13764 25925 13790 25989
rect 13854 25925 13880 25989
rect 13944 25925 13970 25989
rect 14034 25925 14039 25989
rect 13515 25909 14039 25925
rect 13515 25845 13520 25909
rect 13584 25845 13610 25909
rect 13674 25845 13700 25909
rect 13764 25845 13790 25909
rect 13854 25845 13880 25909
rect 13944 25845 13970 25909
rect 14034 25845 14039 25909
rect 13515 25829 14039 25845
rect 13515 25765 13520 25829
rect 13584 25765 13610 25829
rect 13674 25765 13700 25829
rect 13764 25765 13790 25829
rect 13854 25765 13880 25829
rect 13944 25765 13970 25829
rect 14034 25765 14039 25829
rect 13515 25749 14039 25765
rect 13515 25685 13520 25749
rect 13584 25685 13610 25749
rect 13674 25685 13700 25749
rect 13764 25685 13790 25749
rect 13854 25685 13880 25749
rect 13944 25685 13970 25749
rect 14034 25685 14039 25749
rect 13515 25669 14039 25685
rect 13515 25605 13520 25669
rect 13584 25605 13610 25669
rect 13674 25605 13700 25669
rect 13764 25605 13790 25669
rect 13854 25605 13880 25669
rect 13944 25605 13970 25669
rect 14034 25605 14039 25669
rect 13515 25589 14039 25605
rect 13515 25525 13520 25589
rect 13584 25525 13610 25589
rect 13674 25525 13700 25589
rect 13764 25525 13790 25589
rect 13854 25525 13880 25589
rect 13944 25525 13970 25589
rect 14034 25525 14039 25589
rect 13515 25509 14039 25525
rect 13515 25445 13520 25509
rect 13584 25445 13610 25509
rect 13674 25445 13700 25509
rect 13764 25445 13790 25509
rect 13854 25445 13880 25509
rect 13944 25445 13970 25509
rect 14034 25445 14039 25509
rect 13515 25429 14039 25445
rect 13515 25365 13520 25429
rect 13584 25365 13610 25429
rect 13674 25365 13700 25429
rect 13764 25365 13790 25429
rect 13854 25365 13880 25429
rect 13944 25365 13970 25429
rect 14034 25365 14039 25429
rect 13515 25349 14039 25365
rect 13515 25285 13520 25349
rect 13584 25285 13610 25349
rect 13674 25285 13700 25349
rect 13764 25285 13790 25349
rect 13854 25285 13880 25349
rect 13944 25285 13970 25349
rect 14034 25285 14039 25349
rect 13515 25269 14039 25285
rect 13515 25205 13520 25269
rect 13584 25205 13610 25269
rect 13674 25205 13700 25269
rect 13764 25205 13790 25269
rect 13854 25205 13880 25269
rect 13944 25205 13970 25269
rect 14034 25205 14039 25269
rect 13515 25189 14039 25205
rect 13515 25125 13520 25189
rect 13584 25125 13610 25189
rect 13674 25125 13700 25189
rect 13764 25125 13790 25189
rect 13854 25125 13880 25189
rect 13944 25125 13970 25189
rect 14034 25125 14039 25189
rect 13515 25109 14039 25125
rect 13515 25045 13520 25109
rect 13584 25045 13610 25109
rect 13674 25045 13700 25109
rect 13764 25045 13790 25109
rect 13854 25045 13880 25109
rect 13944 25045 13970 25109
rect 14034 25045 14039 25109
rect 13515 25029 14039 25045
rect 13515 24965 13520 25029
rect 13584 24965 13610 25029
rect 13674 24965 13700 25029
rect 13764 24965 13790 25029
rect 13854 24965 13880 25029
rect 13944 24965 13970 25029
rect 14034 24965 14039 25029
rect 13515 24949 14039 24965
rect 13515 24885 13520 24949
rect 13584 24885 13610 24949
rect 13674 24885 13700 24949
rect 13764 24885 13790 24949
rect 13854 24885 13880 24949
rect 13944 24885 13970 24949
rect 14034 24885 14039 24949
rect 13515 24869 14039 24885
rect 13515 24805 13520 24869
rect 13584 24805 13610 24869
rect 13674 24805 13700 24869
rect 13764 24805 13790 24869
rect 13854 24805 13880 24869
rect 13944 24805 13970 24869
rect 14034 24805 14039 24869
rect 13515 24789 14039 24805
rect 13515 24725 13520 24789
rect 13584 24725 13610 24789
rect 13674 24725 13700 24789
rect 13764 24725 13790 24789
rect 13854 24725 13880 24789
rect 13944 24725 13970 24789
rect 14034 24725 14039 24789
rect 13515 24709 14039 24725
rect 13515 24645 13520 24709
rect 13584 24645 13610 24709
rect 13674 24645 13700 24709
rect 13764 24645 13790 24709
rect 13854 24645 13880 24709
rect 13944 24645 13970 24709
rect 14034 24645 14039 24709
rect 13515 24629 14039 24645
rect 13515 24565 13520 24629
rect 13584 24565 13610 24629
rect 13674 24565 13700 24629
rect 13764 24565 13790 24629
rect 13854 24565 13880 24629
rect 13944 24565 13970 24629
rect 14034 24565 14039 24629
rect 13515 24549 14039 24565
rect 13515 24485 13520 24549
rect 13584 24485 13610 24549
rect 13674 24485 13700 24549
rect 13764 24485 13790 24549
rect 13854 24485 13880 24549
rect 13944 24485 13970 24549
rect 14034 24485 14039 24549
rect 13515 24469 14039 24485
rect 13515 24405 13520 24469
rect 13584 24405 13610 24469
rect 13674 24405 13700 24469
rect 13764 24405 13790 24469
rect 13854 24405 13880 24469
rect 13944 24405 13970 24469
rect 14034 24405 14039 24469
rect 13515 24389 14039 24405
rect 13515 24325 13520 24389
rect 13584 24325 13610 24389
rect 13674 24325 13700 24389
rect 13764 24325 13790 24389
rect 13854 24325 13880 24389
rect 13944 24325 13970 24389
rect 14034 24325 14039 24389
rect 13515 24309 14039 24325
rect 13515 24245 13520 24309
rect 13584 24245 13610 24309
rect 13674 24245 13700 24309
rect 13764 24245 13790 24309
rect 13854 24245 13880 24309
rect 13944 24245 13970 24309
rect 14034 24245 14039 24309
rect 13515 24229 14039 24245
rect 13515 24165 13520 24229
rect 13584 24165 13610 24229
rect 13674 24165 13700 24229
rect 13764 24165 13790 24229
rect 13854 24165 13880 24229
rect 13944 24165 13970 24229
rect 14034 24165 14039 24229
rect 13515 24149 14039 24165
rect 13515 24085 13520 24149
rect 13584 24085 13610 24149
rect 13674 24085 13700 24149
rect 13764 24085 13790 24149
rect 13854 24085 13880 24149
rect 13944 24085 13970 24149
rect 14034 24085 14039 24149
rect 13515 24069 14039 24085
rect 13515 24005 13520 24069
rect 13584 24005 13610 24069
rect 13674 24005 13700 24069
rect 13764 24005 13790 24069
rect 13854 24005 13880 24069
rect 13944 24005 13970 24069
rect 14034 24005 14039 24069
rect 13515 23989 14039 24005
rect 13515 23925 13520 23989
rect 13584 23925 13610 23989
rect 13674 23925 13700 23989
rect 13764 23925 13790 23989
rect 13854 23925 13880 23989
rect 13944 23925 13970 23989
rect 14034 23925 14039 23989
rect 13515 23909 14039 23925
rect 13515 23845 13520 23909
rect 13584 23845 13610 23909
rect 13674 23845 13700 23909
rect 13764 23845 13790 23909
rect 13854 23845 13880 23909
rect 13944 23845 13970 23909
rect 14034 23845 14039 23909
rect 13515 23829 14039 23845
rect 13515 23765 13520 23829
rect 13584 23765 13610 23829
rect 13674 23765 13700 23829
rect 13764 23765 13790 23829
rect 13854 23765 13880 23829
rect 13944 23765 13970 23829
rect 14034 23765 14039 23829
rect 13515 23749 14039 23765
rect 13515 23685 13520 23749
rect 13584 23685 13610 23749
rect 13674 23685 13700 23749
rect 13764 23685 13790 23749
rect 13854 23685 13880 23749
rect 13944 23685 13970 23749
rect 14034 23685 14039 23749
rect 13515 23669 14039 23685
rect 13515 23605 13520 23669
rect 13584 23605 13610 23669
rect 13674 23605 13700 23669
rect 13764 23605 13790 23669
rect 13854 23605 13880 23669
rect 13944 23605 13970 23669
rect 14034 23605 14039 23669
rect 13515 23589 14039 23605
rect 13515 23525 13520 23589
rect 13584 23525 13610 23589
rect 13674 23525 13700 23589
rect 13764 23525 13790 23589
rect 13854 23525 13880 23589
rect 13944 23525 13970 23589
rect 14034 23525 14039 23589
rect 13515 23509 14039 23525
rect 13515 23445 13520 23509
rect 13584 23445 13610 23509
rect 13674 23445 13700 23509
rect 13764 23445 13790 23509
rect 13854 23445 13880 23509
rect 13944 23445 13970 23509
rect 14034 23445 14039 23509
rect 13515 23429 14039 23445
rect 13515 23365 13520 23429
rect 13584 23365 13610 23429
rect 13674 23365 13700 23429
rect 13764 23365 13790 23429
rect 13854 23365 13880 23429
rect 13944 23365 13970 23429
rect 14034 23365 14039 23429
rect 13515 23349 14039 23365
rect 13515 23285 13520 23349
rect 13584 23285 13610 23349
rect 13674 23285 13700 23349
rect 13764 23285 13790 23349
rect 13854 23285 13880 23349
rect 13944 23285 13970 23349
rect 14034 23285 14039 23349
rect 13515 23268 14039 23285
rect 13515 23204 13520 23268
rect 13584 23204 13610 23268
rect 13674 23204 13700 23268
rect 13764 23204 13790 23268
rect 13854 23204 13880 23268
rect 13944 23204 13970 23268
rect 14034 23204 14039 23268
rect 13515 23187 14039 23204
rect 13515 23123 13520 23187
rect 13584 23123 13610 23187
rect 13674 23123 13700 23187
rect 13764 23123 13790 23187
rect 13854 23123 13880 23187
rect 13944 23123 13970 23187
rect 14034 23123 14039 23187
rect 13515 23106 14039 23123
rect 13515 23042 13520 23106
rect 13584 23042 13610 23106
rect 13674 23042 13700 23106
rect 13764 23042 13790 23106
rect 13854 23042 13880 23106
rect 13944 23042 13970 23106
rect 14034 23042 14039 23106
rect 13515 23025 14039 23042
rect 13515 22961 13520 23025
rect 13584 22961 13610 23025
rect 13674 22961 13700 23025
rect 13764 22961 13790 23025
rect 13854 22961 13880 23025
rect 13944 22961 13970 23025
rect 14034 22961 14039 23025
rect 13515 22944 14039 22961
rect 13515 22880 13520 22944
rect 13584 22880 13610 22944
rect 13674 22880 13700 22944
rect 13764 22880 13790 22944
rect 13854 22880 13880 22944
rect 13944 22880 13970 22944
rect 14034 22880 14039 22944
rect 13515 22863 14039 22880
rect 13515 22799 13520 22863
rect 13584 22799 13610 22863
rect 13674 22799 13700 22863
rect 13764 22799 13790 22863
rect 13854 22799 13880 22863
rect 13944 22799 13970 22863
rect 14034 22799 14039 22863
rect 13515 22782 14039 22799
rect 13515 22718 13520 22782
rect 13584 22718 13610 22782
rect 13674 22718 13700 22782
rect 13764 22718 13790 22782
rect 13854 22718 13880 22782
rect 13944 22718 13970 22782
rect 14034 22718 14039 22782
rect 13515 22701 14039 22718
rect 13515 22637 13520 22701
rect 13584 22637 13610 22701
rect 13674 22637 13700 22701
rect 13764 22637 13790 22701
rect 13854 22637 13880 22701
rect 13944 22637 13970 22701
rect 14034 22637 14039 22701
rect 13515 22620 14039 22637
rect 13515 22556 13520 22620
rect 13584 22556 13610 22620
rect 13674 22556 13700 22620
rect 13764 22556 13790 22620
rect 13854 22556 13880 22620
rect 13944 22556 13970 22620
rect 14034 22556 14039 22620
rect 13515 22539 14039 22556
rect 13515 22475 13520 22539
rect 13584 22475 13610 22539
rect 13674 22475 13700 22539
rect 13764 22475 13790 22539
rect 13854 22475 13880 22539
rect 13944 22475 13970 22539
rect 14034 22475 14039 22539
rect 13515 22458 14039 22475
rect 13515 22394 13520 22458
rect 13584 22394 13610 22458
rect 13674 22394 13700 22458
rect 13764 22394 13790 22458
rect 13854 22394 13880 22458
rect 13944 22394 13970 22458
rect 14034 22394 14039 22458
rect 13515 22377 14039 22394
rect 13515 22313 13520 22377
rect 13584 22313 13610 22377
rect 13674 22313 13700 22377
rect 13764 22313 13790 22377
rect 13854 22313 13880 22377
rect 13944 22313 13970 22377
rect 14034 22313 14039 22377
rect 13515 22296 14039 22313
rect 13515 22232 13520 22296
rect 13584 22232 13610 22296
rect 13674 22232 13700 22296
rect 13764 22232 13790 22296
rect 13854 22232 13880 22296
rect 13944 22232 13970 22296
rect 14034 22232 14039 22296
rect 13515 22215 14039 22232
rect 13515 22151 13520 22215
rect 13584 22151 13610 22215
rect 13674 22151 13700 22215
rect 13764 22151 13790 22215
rect 13854 22151 13880 22215
rect 13944 22151 13970 22215
rect 14034 22151 14039 22215
rect 13515 22134 14039 22151
rect 13515 22070 13520 22134
rect 13584 22070 13610 22134
rect 13674 22070 13700 22134
rect 13764 22070 13790 22134
rect 13854 22070 13880 22134
rect 13944 22070 13970 22134
rect 14034 22070 14039 22134
rect 13515 22053 14039 22070
rect 13515 21989 13520 22053
rect 13584 21989 13610 22053
rect 13674 21989 13700 22053
rect 13764 21989 13790 22053
rect 13854 21989 13880 22053
rect 13944 21989 13970 22053
rect 14034 21989 14039 22053
rect 13515 21972 14039 21989
rect 13515 21908 13520 21972
rect 13584 21908 13610 21972
rect 13674 21908 13700 21972
rect 13764 21908 13790 21972
rect 13854 21908 13880 21972
rect 13944 21908 13970 21972
rect 14034 21908 14039 21972
rect 13515 21891 14039 21908
rect 13515 21827 13520 21891
rect 13584 21827 13610 21891
rect 13674 21827 13700 21891
rect 13764 21827 13790 21891
rect 13854 21827 13880 21891
rect 13944 21827 13970 21891
rect 14034 21827 14039 21891
rect 13515 21810 14039 21827
rect 13515 21746 13520 21810
rect 13584 21746 13610 21810
rect 13674 21746 13700 21810
rect 13764 21746 13790 21810
rect 13854 21746 13880 21810
rect 13944 21746 13970 21810
rect 14034 21746 14039 21810
rect 13515 21729 14039 21746
rect 13515 21665 13520 21729
rect 13584 21665 13610 21729
rect 13674 21665 13700 21729
rect 13764 21665 13790 21729
rect 13854 21665 13880 21729
rect 13944 21665 13970 21729
rect 14034 21665 14039 21729
rect 13515 21648 14039 21665
rect 13515 21584 13520 21648
rect 13584 21584 13610 21648
rect 13674 21584 13700 21648
rect 13764 21584 13790 21648
rect 13854 21584 13880 21648
rect 13944 21584 13970 21648
rect 14034 21584 14039 21648
rect 13515 21567 14039 21584
rect 13515 21503 13520 21567
rect 13584 21503 13610 21567
rect 13674 21503 13700 21567
rect 13764 21503 13790 21567
rect 13854 21503 13880 21567
rect 13944 21503 13970 21567
rect 14034 21503 14039 21567
rect 13515 21486 14039 21503
rect 13515 21422 13520 21486
rect 13584 21422 13610 21486
rect 13674 21422 13700 21486
rect 13764 21422 13790 21486
rect 13854 21422 13880 21486
rect 13944 21422 13970 21486
rect 14034 21422 14039 21486
rect 13515 21405 14039 21422
rect 13515 21341 13520 21405
rect 13584 21341 13610 21405
rect 13674 21341 13700 21405
rect 13764 21341 13790 21405
rect 13854 21341 13880 21405
rect 13944 21341 13970 21405
rect 14034 21341 14039 21405
rect 13515 21324 14039 21341
rect 13515 21260 13520 21324
rect 13584 21260 13610 21324
rect 13674 21260 13700 21324
rect 13764 21260 13790 21324
rect 13854 21260 13880 21324
rect 13944 21260 13970 21324
rect 14034 21260 14039 21324
rect 13515 21243 14039 21260
rect 13515 21179 13520 21243
rect 13584 21179 13610 21243
rect 13674 21179 13700 21243
rect 13764 21179 13790 21243
rect 13854 21179 13880 21243
rect 13944 21179 13970 21243
rect 14034 21179 14039 21243
rect 13515 21162 14039 21179
rect 13515 21098 13520 21162
rect 13584 21098 13610 21162
rect 13674 21098 13700 21162
rect 13764 21098 13790 21162
rect 13854 21098 13880 21162
rect 13944 21098 13970 21162
rect 14034 21098 14039 21162
rect 13515 21081 14039 21098
rect 13515 21017 13520 21081
rect 13584 21017 13610 21081
rect 13674 21017 13700 21081
rect 13764 21017 13790 21081
rect 13854 21017 13880 21081
rect 13944 21017 13970 21081
rect 14034 21017 14039 21081
rect 13515 21000 14039 21017
rect 13515 20972 13520 21000
rect 1496 20939 1596 20972
rect 1496 20936 1531 20939
rect 977 20919 1531 20936
rect 977 20855 982 20919
rect 1046 20855 1072 20919
rect 1136 20855 1162 20919
rect 1226 20855 1252 20919
rect 1316 20855 1342 20919
rect 1406 20855 1432 20919
rect 1496 20875 1531 20919
rect 1595 20875 1596 20939
rect 1496 20855 1596 20875
rect 977 20854 1596 20855
rect 1471 20842 1596 20854
rect 13420 20939 13520 20972
rect 13420 20875 13421 20939
rect 13485 20936 13520 20939
rect 13584 20936 13610 21000
rect 13674 20936 13700 21000
rect 13764 20936 13790 21000
rect 13854 20936 13880 21000
rect 13944 20936 13970 21000
rect 14034 20936 14039 21000
rect 13485 20919 14039 20936
rect 13485 20875 13520 20919
rect 13420 20855 13520 20875
rect 13584 20855 13610 20919
rect 13674 20855 13700 20919
rect 13764 20855 13790 20919
rect 13854 20855 13880 20919
rect 13944 20855 13970 20919
rect 14034 20855 14039 20919
rect 13420 20854 14039 20855
rect 13420 20842 13545 20854
rect 1311 20825 1736 20827
rect 1140 20783 1265 20816
rect 1140 20719 1141 20783
rect 1205 20719 1265 20783
rect 1140 20686 1265 20719
rect 1311 20761 1312 20825
rect 1376 20761 1401 20825
rect 1465 20761 1491 20825
rect 1555 20761 1581 20825
rect 1645 20761 1671 20825
rect 1735 20761 1736 20825
rect 1311 20709 1736 20761
rect 1311 20645 1312 20709
rect 1376 20645 1401 20709
rect 1465 20645 1491 20709
rect 1555 20645 1581 20709
rect 1645 20645 1671 20709
rect 1735 20645 1736 20709
rect 13280 20825 13705 20827
rect 13280 20761 13281 20825
rect 13345 20761 13371 20825
rect 13435 20761 13461 20825
rect 13525 20761 13551 20825
rect 13615 20761 13640 20825
rect 13704 20761 13705 20825
rect 13280 20709 13705 20761
rect 1311 20593 1736 20645
rect 1311 20529 1312 20593
rect 1376 20529 1401 20593
rect 1465 20529 1491 20593
rect 1555 20529 1581 20593
rect 1645 20529 1671 20593
rect 1735 20529 1736 20593
rect 1752 20631 1877 20664
rect 1752 20567 1812 20631
rect 1876 20567 1877 20631
rect 1752 20534 1877 20567
rect 13139 20631 13264 20664
rect 13139 20567 13140 20631
rect 13204 20567 13264 20631
rect 13139 20534 13264 20567
rect 13280 20645 13281 20709
rect 13345 20645 13371 20709
rect 13435 20645 13461 20709
rect 13525 20645 13551 20709
rect 13615 20645 13640 20709
rect 13704 20645 13705 20709
rect 13719 20823 13843 20824
rect 13719 20759 13749 20823
rect 13813 20759 13843 20823
rect 13719 20712 13843 20759
rect 13849 20816 13916 20849
rect 13849 20752 13851 20816
rect 13915 20752 13916 20816
rect 13849 20719 13916 20752
rect 13719 20648 13749 20712
rect 13813 20648 13843 20712
rect 13719 20647 13843 20648
rect 13280 20593 13705 20645
rect 1311 20527 1736 20529
rect 13280 20529 13281 20593
rect 13345 20529 13371 20593
rect 13435 20529 13461 20593
rect 13525 20529 13551 20593
rect 13615 20529 13640 20593
rect 13704 20529 13705 20593
rect 13280 20527 13705 20529
rect 1631 20505 2056 20507
rect 1464 20469 1589 20502
rect 1464 20405 1524 20469
rect 1588 20405 1589 20469
rect 1464 20372 1589 20405
rect 1631 20441 1632 20505
rect 1696 20441 1721 20505
rect 1785 20441 1811 20505
rect 1875 20441 1901 20505
rect 1965 20441 1991 20505
rect 2055 20441 2056 20505
rect 1631 20389 2056 20441
rect 1631 20325 1632 20389
rect 1696 20325 1721 20389
rect 1785 20325 1811 20389
rect 1875 20325 1901 20389
rect 1965 20325 1991 20389
rect 2055 20325 2056 20389
rect 12960 20505 13385 20507
rect 12960 20441 12961 20505
rect 13025 20441 13051 20505
rect 13115 20441 13141 20505
rect 13205 20441 13231 20505
rect 13295 20441 13320 20505
rect 13384 20441 13385 20505
rect 12960 20389 13385 20441
rect 1631 20273 2056 20325
rect 1631 20209 1632 20273
rect 1696 20209 1721 20273
rect 1785 20209 1811 20273
rect 1875 20209 1901 20273
rect 1965 20209 1991 20273
rect 2055 20209 2056 20273
rect 2077 20306 2202 20339
rect 2077 20242 2137 20306
rect 2201 20242 2202 20306
rect 2077 20209 2202 20242
rect 12814 20306 12939 20339
rect 12814 20242 12815 20306
rect 12879 20242 12939 20306
rect 12814 20209 12939 20242
rect 12960 20325 12961 20389
rect 13025 20325 13051 20389
rect 13115 20325 13141 20389
rect 13205 20325 13231 20389
rect 13295 20325 13320 20389
rect 13384 20325 13385 20389
rect 13427 20469 13552 20502
rect 13427 20405 13428 20469
rect 13492 20405 13552 20469
rect 13427 20372 13552 20405
rect 12960 20273 13385 20325
rect 12960 20209 12961 20273
rect 13025 20209 13051 20273
rect 13115 20209 13141 20273
rect 13205 20209 13231 20273
rect 13295 20209 13320 20273
rect 13384 20209 13385 20273
rect 1631 20207 2056 20209
rect 12960 20207 13385 20209
rect 1955 20181 2380 20183
rect 1792 20141 1917 20174
rect 1792 20077 1852 20141
rect 1916 20077 1917 20141
rect 1792 20044 1917 20077
rect 1955 20117 1956 20181
rect 2020 20117 2045 20181
rect 2109 20117 2135 20181
rect 2199 20117 2225 20181
rect 2289 20117 2315 20181
rect 2379 20117 2380 20181
rect 1955 20065 2380 20117
rect 12636 20181 13061 20183
rect 12636 20117 12637 20181
rect 12701 20117 12727 20181
rect 12791 20117 12817 20181
rect 12881 20117 12907 20181
rect 12971 20117 12996 20181
rect 13060 20117 13061 20181
rect 1955 20001 1956 20065
rect 2020 20001 2045 20065
rect 2109 20001 2135 20065
rect 2199 20001 2225 20065
rect 2289 20001 2315 20065
rect 2379 20001 2380 20065
rect 1955 19949 2380 20001
rect 1955 19885 1956 19949
rect 2020 19885 2045 19949
rect 2109 19885 2135 19949
rect 2199 19885 2225 19949
rect 2289 19885 2315 19949
rect 2379 19885 2380 19949
rect 2455 20070 2867 20071
rect 2455 20006 2456 20070
rect 2520 20006 2571 20070
rect 2635 20006 2686 20070
rect 2750 20006 2802 20070
rect 2866 20006 2867 20070
rect 2455 19950 2867 20006
rect 12149 20070 12561 20071
rect 12149 20006 12150 20070
rect 12214 20006 12266 20070
rect 12330 20006 12381 20070
rect 12445 20006 12496 20070
rect 12560 20006 12561 20070
rect 2455 19886 2456 19950
rect 2520 19886 2571 19950
rect 2635 19886 2686 19950
rect 2750 19886 2802 19950
rect 2866 19886 2867 19950
rect 2455 19885 2867 19886
rect 2881 19955 2971 19988
rect 2881 19891 2906 19955
rect 2970 19891 2971 19955
rect 1955 19883 2380 19885
rect 2881 19858 2971 19891
rect 12045 19955 12135 19988
rect 12045 19891 12046 19955
rect 12110 19891 12135 19955
rect 12045 19858 12135 19891
rect 12149 19950 12561 20006
rect 12149 19886 12150 19950
rect 12214 19886 12266 19950
rect 12330 19886 12381 19950
rect 12445 19886 12496 19950
rect 12560 19886 12561 19950
rect 12149 19885 12561 19886
rect 12636 20065 13061 20117
rect 12636 20001 12637 20065
rect 12701 20001 12727 20065
rect 12791 20001 12817 20065
rect 12881 20001 12907 20065
rect 12971 20001 12996 20065
rect 13060 20001 13061 20065
rect 13099 20141 13224 20174
rect 13099 20077 13100 20141
rect 13164 20077 13224 20141
rect 13099 20044 13224 20077
rect 12636 19949 13061 20001
rect 12636 19885 12637 19949
rect 12701 19885 12727 19949
rect 12791 19885 12817 19949
rect 12881 19885 12907 19949
rect 12971 19885 12996 19949
rect 13060 19885 13061 19949
rect 12636 19883 13061 19885
rect 2292 19844 3114 19846
rect 2133 19800 2258 19833
rect 2133 19736 2193 19800
rect 2257 19736 2258 19800
rect 2133 19703 2258 19736
rect 2292 19780 2293 19844
rect 2357 19780 2377 19844
rect 2441 19780 2461 19844
rect 2525 19780 2545 19844
rect 2609 19780 2629 19844
rect 2693 19780 2713 19844
rect 2777 19780 2797 19844
rect 2861 19780 2881 19844
rect 2945 19780 2965 19844
rect 3029 19780 3049 19844
rect 3113 19780 3114 19844
rect 2292 19728 3114 19780
rect 2292 19664 2293 19728
rect 2357 19664 2377 19728
rect 2441 19664 2461 19728
rect 2525 19664 2545 19728
rect 2609 19664 2629 19728
rect 2693 19664 2713 19728
rect 2777 19664 2797 19728
rect 2861 19664 2881 19728
rect 2945 19664 2965 19728
rect 3029 19664 3049 19728
rect 3113 19664 3114 19728
rect 11902 19844 12724 19846
rect 11902 19780 11903 19844
rect 11967 19780 11987 19844
rect 12051 19780 12071 19844
rect 12135 19780 12155 19844
rect 12219 19780 12239 19844
rect 12303 19780 12323 19844
rect 12387 19780 12407 19844
rect 12471 19780 12491 19844
rect 12555 19780 12575 19844
rect 12639 19780 12659 19844
rect 12723 19780 12724 19844
rect 11902 19728 12724 19780
rect 2292 19612 3114 19664
rect 2292 19548 2293 19612
rect 2357 19548 2377 19612
rect 2441 19548 2461 19612
rect 2525 19548 2545 19612
rect 2609 19548 2629 19612
rect 2693 19548 2713 19612
rect 2777 19548 2797 19612
rect 2861 19548 2881 19612
rect 2945 19548 2965 19612
rect 3029 19548 3049 19612
rect 3113 19548 3114 19612
rect 3123 19707 3247 19708
rect 3123 19643 3153 19707
rect 3217 19643 3247 19707
rect 3123 19614 3247 19643
rect 3123 19550 3153 19614
rect 3217 19550 3247 19614
rect 3123 19549 3247 19550
rect 11769 19707 11893 19708
rect 11769 19643 11799 19707
rect 11863 19643 11893 19707
rect 11769 19614 11893 19643
rect 11769 19550 11799 19614
rect 11863 19550 11893 19614
rect 11769 19549 11893 19550
rect 11902 19664 11903 19728
rect 11967 19664 11987 19728
rect 12051 19664 12071 19728
rect 12135 19664 12155 19728
rect 12219 19664 12239 19728
rect 12303 19664 12323 19728
rect 12387 19664 12407 19728
rect 12471 19664 12491 19728
rect 12555 19664 12575 19728
rect 12639 19664 12659 19728
rect 12723 19664 12724 19728
rect 12758 19800 12883 19833
rect 12758 19736 12759 19800
rect 12823 19736 12883 19800
rect 12758 19703 12883 19736
rect 11902 19612 12724 19664
rect 2292 19546 3114 19548
rect 11902 19548 11903 19612
rect 11967 19548 11987 19612
rect 12051 19548 12071 19612
rect 12135 19548 12155 19612
rect 12219 19548 12239 19612
rect 12303 19548 12323 19612
rect 12387 19548 12407 19612
rect 12471 19548 12491 19612
rect 12555 19548 12575 19612
rect 12639 19548 12659 19612
rect 12723 19548 12724 19612
rect 11902 19546 12724 19548
rect 3916 7963 5155 8038
rect 3916 7419 3977 7963
rect 5081 7419 5155 7963
rect 3916 7348 5155 7419
rect 9753 7965 10992 8038
rect 9753 7421 9820 7965
rect 10924 7421 10992 7965
rect 9753 7348 10992 7421
rect 2423 6025 3607 6053
rect 2423 5213 3607 5241
rect 11297 6024 12481 6052
rect 11297 5212 12481 5240
rect 858 3611 2098 3678
rect 858 3067 924 3611
rect 2028 3067 2098 3611
rect 858 2999 2098 3067
rect 12858 3643 14098 3678
rect 12858 3019 12928 3643
rect 14032 3019 14098 3643
rect 12858 2991 14098 3019
use sky130_fd_io__com_busses_esd  sky130_fd_io__com_busses_esd_0
timestamp 1688980957
transform 1 0 8 0 1 550
box 0 -142 15000 39451
<< properties >>
string GDS_END 5216472
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 4497834
<< end >>
