magic
tech sky130B
magscale 1 2
timestamp 1688980957
use sky130_fd_pr__dfl1sd__example_5595914180815  sky130_fd_pr__dfl1sd__example_5595914180815_0
timestamp 1688980957
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_0
timestamp 1688980957
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_0
timestamp 1688980957
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 48384088
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48382646
<< end >>
