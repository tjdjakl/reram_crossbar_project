magic
tech sky130B
magscale 1 2
timestamp 1700640585
<< metal1 >>
rect 31506 22890 31706 23090
rect 33370 22920 33380 23080
rect 33560 22920 33570 23080
rect 31412 22498 31612 22698
rect 31400 21852 31600 22052
rect 31412 21386 31612 21586
rect 31504 21056 31704 21256
rect 33370 21040 33380 21180
rect 33560 21040 33570 21180
rect 34114 20681 34124 20821
rect 34282 20681 34292 20821
rect 38090 20720 38100 20880
rect 38260 20720 38270 20880
rect 33160 19620 34040 19820
rect 38664 19646 38864 19846
rect 35070 18860 35080 19000
rect 35240 18860 35250 19000
rect 34112 18491 34122 18631
rect 34280 18491 34290 18631
rect 38090 18520 38100 18680
rect 38260 18520 38270 18680
rect 33160 17420 34000 17620
rect 38664 17446 38864 17646
rect 35070 16660 35080 16800
rect 35240 16660 35250 16800
rect 34114 16306 34124 16446
rect 34282 16306 34292 16446
rect 38090 16340 38100 16500
rect 38260 16340 38270 16500
rect 33160 15220 34000 15420
rect 38664 15246 38864 15446
rect 35070 14440 35080 14580
rect 35240 14440 35250 14580
rect 34112 14092 34122 14232
rect 34280 14092 34290 14232
rect 38090 14120 38100 14280
rect 38260 14120 38270 14280
rect 33160 13020 34000 13220
rect 38664 13046 38864 13246
rect 35070 12260 35080 12400
rect 35240 12260 35250 12400
rect 34115 11900 34125 12040
rect 34283 11900 34293 12040
rect 38090 11920 38100 12080
rect 38260 11920 38270 12080
rect 33160 10820 34000 11020
rect 38664 10846 38864 11046
rect 35070 10040 35080 10180
rect 35240 10040 35250 10180
rect 34115 9696 34125 9836
rect 34283 9696 34293 9836
rect 38090 9720 38100 9880
rect 38260 9720 38270 9880
rect 33160 8620 34000 8820
rect 38664 8646 38864 8846
rect 35070 7840 35080 7980
rect 35240 7840 35250 7980
rect 34115 7491 34125 7631
rect 34283 7491 34293 7631
rect 38090 7520 38100 7680
rect 38260 7520 38270 7680
rect 33160 6420 34000 6620
rect 38664 6446 38864 6646
rect 35070 5640 35080 5780
rect 35240 5640 35250 5780
rect 34112 5297 34122 5437
rect 34280 5297 34290 5437
rect 38090 5320 38100 5480
rect 38260 5320 38270 5480
rect 33160 4220 34000 4420
rect 38664 4246 38864 4446
rect 35070 3440 35080 3580
rect 35240 3440 35250 3580
<< via1 >>
rect 33380 22920 33560 23080
rect 33380 21040 33560 21180
rect 34124 20681 34282 20821
rect 38100 20720 38260 20880
rect 35080 18860 35240 19000
rect 34122 18491 34280 18631
rect 38100 18520 38260 18680
rect 35080 16660 35240 16800
rect 34124 16306 34282 16446
rect 38100 16340 38260 16500
rect 35080 14440 35240 14580
rect 34122 14092 34280 14232
rect 38100 14120 38260 14280
rect 35080 12260 35240 12400
rect 34125 11900 34283 12040
rect 38100 11920 38260 12080
rect 35080 10040 35240 10180
rect 34125 9696 34283 9836
rect 38100 9720 38260 9880
rect 35080 7840 35240 7980
rect 34125 7491 34283 7631
rect 38100 7520 38260 7680
rect 35080 5640 35240 5780
rect 34122 5297 34280 5437
rect 38100 5320 38260 5480
rect 35080 3440 35240 3580
<< metal2 >>
rect 33380 23080 33560 23090
rect 33380 22910 33560 22920
rect 33986 21997 34133 22007
rect 33986 21870 34133 21880
rect 33380 21180 33560 21190
rect 33380 21030 33560 21040
rect 38100 20880 38260 20890
rect 34124 20821 34282 20831
rect 38100 20710 38260 20720
rect 34124 20671 34282 20681
rect 33160 20180 33360 20240
rect 33720 20180 33840 20190
rect 33160 20060 33720 20180
rect 33840 20060 36280 20180
rect 33160 20040 33360 20060
rect 33720 20050 33840 20060
rect 36140 19720 36280 20060
rect 33160 19340 33360 19400
rect 33420 19340 33540 19350
rect 33160 19220 33420 19340
rect 33540 19220 36240 19340
rect 33160 19200 33360 19220
rect 33420 19210 33540 19220
rect 35080 19000 35240 19010
rect 35080 18850 35240 18860
rect 38100 18680 38260 18690
rect 34122 18631 34280 18641
rect 38100 18510 38260 18520
rect 34122 18481 34280 18491
rect 33720 17980 33840 17990
rect 33840 17860 36280 17980
rect 33720 17850 33840 17860
rect 36140 17520 36280 17860
rect 33420 17140 33540 17150
rect 33540 17020 36240 17140
rect 33420 17010 33540 17020
rect 35080 16800 35240 16810
rect 35080 16650 35240 16660
rect 38100 16500 38260 16510
rect 34124 16446 34282 16456
rect 38100 16330 38260 16340
rect 34124 16296 34282 16306
rect 33720 15780 33840 15790
rect 33840 15660 36280 15780
rect 33720 15650 33840 15660
rect 36140 15320 36280 15660
rect 33420 14940 33540 14950
rect 33540 14820 36240 14940
rect 33420 14810 33540 14820
rect 35080 14580 35240 14590
rect 35080 14430 35240 14440
rect 38100 14280 38260 14290
rect 34122 14232 34280 14242
rect 38100 14110 38260 14120
rect 34122 14082 34280 14092
rect 33720 13580 33840 13590
rect 33840 13460 36280 13580
rect 33720 13450 33840 13460
rect 36140 13120 36280 13460
rect 33420 12740 33540 12750
rect 33540 12620 36240 12740
rect 33420 12610 33540 12620
rect 35080 12400 35240 12410
rect 35080 12250 35240 12260
rect 38100 12080 38260 12090
rect 34125 12040 34283 12050
rect 38100 11910 38260 11920
rect 34125 11890 34283 11900
rect 33720 11380 33840 11390
rect 33840 11260 36280 11380
rect 33720 11250 33840 11260
rect 36140 10920 36280 11260
rect 33420 10540 33540 10550
rect 33540 10420 36240 10540
rect 33420 10410 33540 10420
rect 35080 10180 35240 10190
rect 35080 10030 35240 10040
rect 38100 9880 38260 9890
rect 34125 9836 34283 9846
rect 38100 9710 38260 9720
rect 34125 9686 34283 9696
rect 33720 9180 33840 9190
rect 33840 9060 36280 9180
rect 33720 9050 33840 9060
rect 36140 8720 36280 9060
rect 33420 8340 33540 8350
rect 33540 8220 36240 8340
rect 33420 8210 33540 8220
rect 35080 7980 35240 7990
rect 35080 7830 35240 7840
rect 38100 7680 38260 7690
rect 34125 7631 34283 7641
rect 38100 7510 38260 7520
rect 34125 7481 34283 7491
rect 33720 6980 33840 6990
rect 33840 6860 36280 6980
rect 33720 6850 33840 6860
rect 36140 6520 36280 6860
rect 33420 6140 33540 6150
rect 33540 6020 36240 6140
rect 33420 6010 33540 6020
rect 35080 5780 35240 5790
rect 35080 5630 35240 5640
rect 38100 5480 38260 5490
rect 34122 5437 34280 5447
rect 38100 5310 38260 5320
rect 34122 5287 34280 5297
rect 33720 4780 33840 4790
rect 33840 4660 36280 4780
rect 33720 4650 33840 4660
rect 36140 4320 36280 4660
rect 33420 3940 33540 3950
rect 33540 3820 36240 3940
rect 33420 3810 33540 3820
rect 35080 3580 35240 3590
rect 35080 3430 35240 3440
<< via2 >>
rect 33380 22920 33560 23080
rect 33986 21880 34133 21997
rect 33380 21040 33560 21180
rect 34124 20681 34282 20821
rect 38100 20720 38260 20880
rect 33720 20060 33840 20180
rect 33420 19220 33540 19340
rect 35080 18860 35240 19000
rect 34122 18491 34280 18631
rect 38100 18520 38260 18680
rect 33720 17860 33840 17980
rect 33420 17020 33540 17140
rect 35080 16660 35240 16800
rect 34124 16306 34282 16446
rect 38100 16340 38260 16500
rect 33720 15660 33840 15780
rect 33420 14820 33540 14940
rect 35080 14440 35240 14580
rect 34122 14092 34280 14232
rect 38100 14120 38260 14280
rect 33720 13460 33840 13580
rect 33420 12620 33540 12740
rect 35080 12260 35240 12400
rect 34125 11900 34283 12040
rect 38100 11920 38260 12080
rect 33720 11260 33840 11380
rect 33420 10420 33540 10540
rect 35080 10040 35240 10180
rect 34125 9696 34283 9836
rect 38100 9720 38260 9880
rect 33720 9060 33840 9180
rect 33420 8220 33540 8340
rect 35080 7840 35240 7980
rect 34125 7491 34283 7631
rect 38100 7520 38260 7680
rect 33720 6860 33840 6980
rect 33420 6020 33540 6140
rect 35080 5640 35240 5780
rect 34122 5297 34280 5437
rect 38100 5320 38260 5480
rect 33720 4660 33840 4780
rect 33420 3820 33540 3940
rect 35080 3440 35240 3580
<< metal3 >>
rect 33370 23080 33570 23085
rect 33370 22920 33380 23080
rect 33560 22940 36240 23080
rect 33560 22920 33570 22940
rect 33370 22915 33570 22920
rect 34124 22002 34282 22007
rect 33976 21997 34282 22002
rect 33976 21880 33986 21997
rect 34133 21880 34282 21997
rect 33976 21875 34282 21880
rect 33370 21180 33570 21185
rect 33370 21040 33380 21180
rect 33560 21040 33570 21180
rect 33370 21035 33570 21040
rect 34124 20826 34282 21875
rect 35070 21040 35080 21160
rect 35240 21040 35250 21160
rect 34114 20821 34292 20826
rect 34114 20681 34124 20821
rect 34282 20681 34292 20821
rect 34114 20676 34292 20681
rect 33710 20180 33850 20185
rect 33710 20060 33720 20180
rect 33840 20060 33850 20180
rect 33710 20055 33850 20060
rect 33410 19340 33550 19345
rect 33410 19220 33420 19340
rect 33540 19220 33550 19340
rect 33410 19215 33550 19220
rect 33420 17145 33540 19215
rect 33720 17985 33840 20055
rect 34124 18636 34280 20676
rect 35080 19005 35240 21040
rect 36100 20880 36240 22940
rect 38090 20880 38270 20885
rect 36100 20720 38100 20880
rect 38260 20720 38500 20880
rect 38090 20715 38270 20720
rect 35070 19000 35250 19005
rect 35070 18860 35080 19000
rect 35240 18860 35250 19000
rect 35070 18855 35250 18860
rect 34112 18631 34290 18636
rect 34112 18491 34122 18631
rect 34280 18491 34290 18631
rect 34112 18486 34290 18491
rect 33710 17980 33850 17985
rect 33710 17860 33720 17980
rect 33840 17860 33850 17980
rect 33710 17855 33850 17860
rect 33410 17140 33550 17145
rect 33410 17020 33420 17140
rect 33540 17020 33550 17140
rect 33410 17015 33550 17020
rect 33420 14945 33540 17015
rect 33720 15785 33840 17855
rect 34124 16451 34280 18486
rect 35080 16805 35240 18855
rect 38090 18680 38270 18685
rect 38340 18680 38480 20720
rect 38090 18520 38100 18680
rect 38260 18520 38480 18680
rect 38090 18515 38270 18520
rect 35070 16800 35250 16805
rect 35070 16660 35080 16800
rect 35240 16660 35250 16800
rect 35070 16655 35250 16660
rect 34114 16446 34292 16451
rect 34114 16306 34124 16446
rect 34282 16306 34292 16446
rect 34114 16301 34292 16306
rect 33710 15780 33850 15785
rect 33710 15660 33720 15780
rect 33840 15660 33850 15780
rect 33710 15655 33850 15660
rect 33410 14940 33550 14945
rect 33410 14820 33420 14940
rect 33540 14820 33550 14940
rect 33410 14815 33550 14820
rect 33420 12745 33540 14815
rect 33720 13585 33840 15655
rect 34124 14237 34280 16301
rect 35080 14585 35240 16655
rect 38090 16500 38270 16505
rect 38340 16500 38480 18520
rect 38090 16340 38100 16500
rect 38260 16340 38480 16500
rect 38090 16335 38270 16340
rect 35070 14580 35250 14585
rect 35070 14440 35080 14580
rect 35240 14440 35250 14580
rect 35070 14435 35250 14440
rect 34112 14232 34290 14237
rect 34112 14092 34122 14232
rect 34280 14092 34290 14232
rect 34112 14087 34290 14092
rect 33710 13580 33850 13585
rect 33710 13460 33720 13580
rect 33840 13460 33850 13580
rect 33710 13455 33850 13460
rect 33410 12740 33550 12745
rect 33410 12620 33420 12740
rect 33540 12620 33550 12740
rect 33410 12615 33550 12620
rect 33420 10545 33540 12615
rect 33720 11385 33840 13455
rect 34124 12045 34280 14087
rect 35080 12405 35240 14435
rect 38090 14280 38270 14285
rect 38340 14280 38480 16340
rect 38090 14120 38100 14280
rect 38260 14120 38480 14280
rect 38090 14115 38270 14120
rect 35070 12400 35250 12405
rect 35070 12260 35080 12400
rect 35240 12260 35250 12400
rect 35070 12255 35250 12260
rect 34115 12040 34293 12045
rect 34115 11900 34125 12040
rect 34283 11900 34293 12040
rect 34115 11895 34293 11900
rect 33710 11380 33850 11385
rect 33710 11260 33720 11380
rect 33840 11260 33850 11380
rect 33710 11255 33850 11260
rect 33410 10540 33550 10545
rect 33410 10420 33420 10540
rect 33540 10420 33550 10540
rect 33410 10415 33550 10420
rect 33420 8345 33540 10415
rect 33720 9185 33840 11255
rect 34124 9841 34280 11895
rect 35080 10185 35240 12255
rect 38090 12080 38270 12085
rect 38340 12080 38480 14120
rect 38090 11920 38100 12080
rect 38260 11920 38480 12080
rect 38090 11915 38270 11920
rect 35070 10180 35250 10185
rect 35070 10040 35080 10180
rect 35240 10040 35250 10180
rect 35070 10035 35250 10040
rect 34115 9836 34293 9841
rect 34115 9696 34125 9836
rect 34283 9696 34293 9836
rect 34115 9691 34293 9696
rect 33710 9180 33850 9185
rect 33710 9060 33720 9180
rect 33840 9060 33850 9180
rect 33710 9055 33850 9060
rect 33410 8340 33550 8345
rect 33410 8220 33420 8340
rect 33540 8220 33550 8340
rect 33410 8215 33550 8220
rect 33420 6145 33540 8215
rect 33720 6985 33840 9055
rect 34124 7636 34280 9691
rect 35080 7985 35240 10035
rect 38090 9880 38270 9885
rect 38340 9880 38480 11920
rect 38090 9720 38100 9880
rect 38260 9720 38480 9880
rect 38090 9715 38270 9720
rect 35070 7980 35250 7985
rect 35070 7840 35080 7980
rect 35240 7840 35250 7980
rect 35070 7835 35250 7840
rect 34115 7631 34293 7636
rect 34115 7491 34125 7631
rect 34283 7491 34293 7631
rect 34115 7486 34293 7491
rect 33710 6980 33850 6985
rect 33710 6860 33720 6980
rect 33840 6860 33850 6980
rect 33710 6855 33850 6860
rect 33410 6140 33550 6145
rect 33410 6020 33420 6140
rect 33540 6020 33550 6140
rect 33410 6015 33550 6020
rect 33420 3945 33540 6015
rect 33720 4785 33840 6855
rect 34124 5442 34280 7486
rect 35080 5785 35240 7835
rect 38090 7680 38270 7685
rect 38340 7680 38480 9720
rect 38090 7520 38100 7680
rect 38260 7520 38480 7680
rect 38090 7515 38270 7520
rect 35070 5780 35250 5785
rect 35070 5640 35080 5780
rect 35240 5640 35250 5780
rect 35070 5635 35250 5640
rect 34112 5437 34290 5442
rect 34112 5297 34122 5437
rect 34280 5297 34290 5437
rect 34112 5292 34290 5297
rect 33710 4780 33850 4785
rect 33710 4660 33720 4780
rect 33840 4660 33850 4780
rect 33710 4655 33850 4660
rect 33410 3940 33550 3945
rect 33410 3820 33420 3940
rect 33540 3820 33550 3940
rect 33410 3815 33550 3820
rect 35080 3585 35240 5635
rect 38090 5480 38270 5485
rect 38340 5480 38480 7520
rect 38090 5320 38100 5480
rect 38260 5320 38480 5480
rect 38090 5315 38270 5320
rect 35070 3580 35250 3585
rect 35070 3440 35080 3580
rect 35240 3440 35250 3580
rect 35070 3435 35250 3440
<< via3 >>
rect 33380 21040 33560 21180
rect 35080 21040 35240 21160
<< metal4 >>
rect 33379 21180 33561 21181
rect 33379 21040 33380 21180
rect 33560 21160 33561 21180
rect 35079 21160 35241 21161
rect 33560 21040 35080 21160
rect 35240 21040 35241 21160
rect 33379 21039 33561 21040
rect 35079 21039 35241 21040
use 1LineBitInput  x1
timestamp 1700640585
transform 1 0 29628 0 1 15640
box 4372 3160 9236 5276
use 1LineBitInput  x2
timestamp 1700640585
transform 1 0 29628 0 1 13440
box 4372 3160 9236 5276
use 1LineBitInput  x3
timestamp 1700640585
transform 1 0 29628 0 1 11240
box 4372 3160 9236 5276
use 1LineBitInput  x4
timestamp 1700640585
transform 1 0 29628 0 1 9040
box 4372 3160 9236 5276
use 1LineBitInput  x5
timestamp 1700640585
transform 1 0 29628 0 1 6840
box 4372 3160 9236 5276
use 1LineBitInput  x6
timestamp 1700640585
transform 1 0 29628 0 1 4640
box 4372 3160 9236 5276
use 1LineBitInput  x7
timestamp 1700640585
transform 1 0 29628 0 1 2440
box 4372 3160 9236 5276
use 1LineBitInput  x8
timestamp 1700640585
transform 1 0 29628 0 1 240
box 4372 3160 9236 5276
use 2-1MUX  x9
timestamp 1700640585
transform 1 0 32336 0 1 20400
box -936 600 1824 2716
<< labels >>
flabel metal1 31506 22890 31706 23090 0 FreeSans 256 0 0 0 VDD
port 23 nsew
flabel metal1 31504 21056 31704 21256 0 FreeSans 256 0 0 0 VSS
port 24 nsew
flabel metal1 38664 4246 38864 4446 0 FreeSans 256 0 0 0 BL_IN8
port 22 nsew
flabel metal1 38664 6446 38864 6646 0 FreeSans 256 0 0 0 BL_IN7
port 21 nsew
flabel metal1 38664 8646 38864 8846 0 FreeSans 256 0 0 0 BL_IN6
port 20 nsew
flabel metal1 38664 10846 38864 11046 0 FreeSans 256 0 0 0 BL_IN5
port 19 nsew
flabel metal1 38664 13046 38864 13246 0 FreeSans 256 0 0 0 BL_IN4
port 17 nsew
flabel metal1 38664 15246 38864 15446 0 FreeSans 256 0 0 0 BL_IN3
port 16 nsew
flabel metal1 38664 17446 38864 17646 0 FreeSans 256 0 0 0 BL_IN2
port 15 nsew
flabel metal1 38664 19646 38864 19846 0 FreeSans 256 0 0 0 BL_IN1
port 14 nsew
flabel metal1 31400 21852 31600 22052 0 FreeSans 256 0 0 0 Write_Select
port 0 nsew
flabel metal1 31412 22498 31612 22698 0 FreeSans 256 0 0 0 Write_Voltage
port 1 nsew
flabel metal1 31412 21386 31612 21586 0 FreeSans 256 0 0 0 Form_Voltage
port 2 nsew
flabel metal2 33160 20040 33360 20240 0 FreeSans 256 0 0 0 Write_Form_Select
port 12 nsew
flabel metal2 33160 19200 33360 19400 0 FreeSans 256 0 0 0 MAC_Voltage
port 13 nsew
flabel metal1 33160 19620 33360 19820 0 FreeSans 256 0 0 0 BL_LA_IN1
port 3 nsew
flabel metal1 33160 17420 33360 17620 0 FreeSans 256 0 0 0 BL_LA_IN2
port 11 nsew
flabel metal1 33160 15220 33360 15420 0 FreeSans 256 0 0 0 BL_LA_IN3
port 4 nsew
flabel metal1 33160 13020 33360 13220 0 FreeSans 256 0 0 0 BL_LA_IN4
port 7 nsew
flabel metal1 33160 10820 33360 11020 0 FreeSans 256 0 0 0 BL_LA_IN5
port 8 nsew
flabel metal1 33160 8620 33360 8820 0 FreeSans 256 0 0 0 BL_LA_IN6
port 5 nsew
flabel metal1 33160 6420 33360 6620 0 FreeSans 256 0 0 0 BL_LA_IN7
port 9 nsew
flabel metal1 33160 4220 33360 4420 0 FreeSans 256 0 0 0 BL_LA_IN8
port 10 nsew
<< end >>
