magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 3 157 272 203
rect 3 21 808 157
rect 25 -17 59 21
<< locali >>
rect 105 305 156 493
rect 105 162 139 305
rect 269 199 335 323
rect 369 199 427 275
rect 105 51 156 162
rect 610 271 706 331
rect 654 153 706 271
rect 746 153 798 331
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 37 289 71 527
rect 190 447 256 527
rect 500 474 534 493
rect 308 440 534 474
rect 575 451 641 485
rect 308 395 342 440
rect 190 361 342 395
rect 488 413 534 440
rect 37 17 71 186
rect 190 265 224 361
rect 395 343 429 381
rect 488 379 570 413
rect 173 199 224 265
rect 395 309 502 343
rect 468 165 502 309
rect 323 131 502 165
rect 536 174 570 379
rect 607 401 641 451
rect 675 435 725 527
rect 759 401 793 493
rect 607 367 793 401
rect 536 140 606 174
rect 190 17 276 106
rect 323 51 357 131
rect 391 17 538 97
rect 572 51 606 140
rect 721 17 801 119
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 269 199 335 323 6 A1_N
port 1 nsew signal input
rlabel locali s 369 199 427 275 6 A2_N
port 2 nsew signal input
rlabel locali s 746 153 798 331 6 B1
port 3 nsew signal input
rlabel locali s 654 153 706 271 6 B2
port 4 nsew signal input
rlabel locali s 610 271 706 331 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 25 -17 59 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 3 21 808 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 3 157 272 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 105 51 156 162 6 X
port 9 nsew signal output
rlabel locali s 105 162 139 305 6 X
port 9 nsew signal output
rlabel locali s 105 305 156 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3934450
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3926722
<< end >>
