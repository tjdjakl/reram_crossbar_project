magic
tech sky130B
magscale 1 2
timestamp 1700640585
<< metal1 >>
rect 71478 40048 71678 40248
rect 59149 38559 59350 38759
rect 68568 38646 68768 38846
rect 66314 38273 66514 38473
rect 58808 38019 58818 38180
rect 58980 38019 58990 38180
rect 71478 31048 71678 31248
rect 58810 29020 58820 29181
rect 58982 29020 58992 29181
rect 71478 22048 71678 22248
rect 58810 20020 58820 20181
rect 58982 20020 58992 20181
rect 34080 15572 34280 15772
rect 32180 14776 32380 14976
rect 45188 14728 45388 14928
rect 46052 14708 46252 14908
rect 44610 13680 44620 13840
rect 44780 13680 44790 13840
rect 48596 13342 48796 13542
rect 71478 13048 71678 13248
rect 32180 12576 32380 12776
rect 44610 11480 44620 11640
rect 44780 11480 44790 11640
rect 48596 11142 48796 11342
rect 58810 11020 58820 11181
rect 58982 11020 58992 11181
rect 32180 10376 32380 10576
rect 44610 9280 44620 9440
rect 44780 9280 44790 9440
rect 48596 8942 48796 9142
rect 32180 8176 32380 8376
rect 44610 7080 44620 7240
rect 44780 7080 44790 7240
rect 48596 6742 48796 6942
rect 32180 5976 32380 6176
rect 44610 4880 44620 5040
rect 44780 4880 44790 5040
rect 48596 4542 48796 4742
rect 71478 4048 71678 4248
rect 32180 3776 32380 3976
rect 44610 2680 44620 2840
rect 44780 2680 44790 2840
rect 48596 2342 48796 2542
rect 58810 2020 58820 2181
rect 58982 2020 58992 2181
rect 32180 1576 32380 1776
rect 44610 480 44620 640
rect 44780 480 44790 640
rect 48576 142 48776 342
rect 32180 -624 32380 -424
rect 35230 -1694 35430 -1494
rect 44610 -1720 44620 -1560
rect 44780 -1720 44790 -1560
rect 48160 -1730 48360 -1530
rect 48595 -2058 48796 -1858
rect 30432 -2388 30632 -2188
rect 45186 -2568 45386 -2368
rect 30420 -2856 30620 -2656
rect 30432 -3502 30632 -3302
rect 30392 -4922 30592 -4722
rect 71478 -4952 71678 -4752
rect 30380 -5568 30580 -5368
rect 30392 -6034 30592 -5834
rect 32942 -6742 33142 -6542
rect 58810 -6980 58820 -6819
rect 58982 -6980 58992 -6819
rect 32836 -7780 33036 -7580
rect 34484 -7759 34494 -7619
rect 34654 -7759 34664 -7619
rect 32836 -10180 33036 -9980
rect 34483 -10160 34493 -10020
rect 34653 -10160 34663 -10020
rect 32836 -12580 33036 -12380
rect 34479 -12557 34489 -12417
rect 34649 -12557 34659 -12417
rect 71478 -13952 71678 -13752
rect 32836 -14981 33036 -14780
rect 34483 -14954 34493 -14814
rect 34653 -14954 34663 -14814
rect 58810 -15980 58820 -15819
rect 58982 -15980 58992 -15819
rect 32835 -17380 33035 -17180
rect 34488 -17347 34498 -17207
rect 34658 -17347 34668 -17207
rect 32836 -19780 33036 -19580
rect 34486 -19749 34496 -19609
rect 34656 -19749 34666 -19609
rect 32834 -22180 33036 -21980
rect 34488 -22151 34498 -22011
rect 34658 -22151 34668 -22011
rect 71478 -22952 71678 -22752
rect 32836 -24580 33036 -24380
rect 34490 -24560 34500 -24420
rect 34660 -24560 34670 -24420
rect 58810 -24980 58820 -24819
rect 58982 -24980 58992 -24819
rect 32940 -25376 33140 -25176
<< via1 >>
rect 58818 38019 58980 38180
rect 58820 29020 58982 29181
rect 58820 20020 58982 20181
rect 44620 13680 44780 13840
rect 44620 11480 44780 11640
rect 58820 11020 58982 11181
rect 44620 9280 44780 9440
rect 44620 7080 44780 7240
rect 44620 4880 44780 5040
rect 44620 2680 44780 2840
rect 58820 2020 58982 2181
rect 44620 480 44780 640
rect 44620 -1720 44780 -1560
rect 58820 -6980 58982 -6819
rect 34494 -7759 34654 -7619
rect 34493 -10160 34653 -10020
rect 34489 -12557 34649 -12417
rect 34493 -14954 34653 -14814
rect 58820 -15980 58982 -15819
rect 34498 -17347 34658 -17207
rect 34496 -19749 34656 -19609
rect 34498 -22151 34658 -22011
rect 34500 -24560 34660 -24420
rect 58820 -24980 58982 -24819
<< metal2 >>
rect 58818 38181 58980 38190
rect 52856 38180 58980 38181
rect 51540 38020 58818 38180
rect 51540 18360 51720 38020
rect 58818 38009 58980 38019
rect 58820 29181 58982 29191
rect 52865 29180 58820 29181
rect 38200 18200 51720 18360
rect 51980 29020 58820 29180
rect 37714 14908 37854 14918
rect 37714 14796 37854 14806
rect 38200 13520 38360 18200
rect 51980 18000 52160 29020
rect 58820 29010 58982 29020
rect 58820 20181 58982 20191
rect 52855 20180 58820 20181
rect 38200 13350 38360 13360
rect 38880 17840 52160 18000
rect 52520 20020 58820 20180
rect 37714 12708 37854 12718
rect 37714 12596 37854 12606
rect 38880 11320 39040 17840
rect 52520 17600 52660 20020
rect 58820 20010 58982 20020
rect 38880 11170 39040 11180
rect 39580 17420 52660 17600
rect 37714 10508 37854 10518
rect 37714 10396 37854 10406
rect 39580 9180 39740 17420
rect 39580 9010 39740 9020
rect 40280 16160 40440 16162
rect 40280 16000 52740 16160
rect 37714 8308 37854 8318
rect 37714 8196 37854 8206
rect 40280 7080 40440 16000
rect 44620 13840 44780 13850
rect 44620 13670 44780 13680
rect 44620 11640 44780 11650
rect 44620 11470 44780 11480
rect 52560 11180 52740 16000
rect 58820 11181 58982 11191
rect 52899 11180 58820 11181
rect 52560 11020 58820 11180
rect 58820 11010 58982 11020
rect 44620 9440 44780 9450
rect 44620 9270 44780 9280
rect 44620 7240 44780 7250
rect 44620 7070 44780 7080
rect 40280 6910 40440 6920
rect 37714 6108 37854 6118
rect 37714 5996 37854 6006
rect 44620 5040 44780 5050
rect 44620 4870 44780 4880
rect 37714 3908 37854 3918
rect 37714 3796 37854 3806
rect 44620 2840 44780 2850
rect 44620 2670 44780 2680
rect 58820 2181 58982 2191
rect 52899 2180 58820 2181
rect 52620 2020 58820 2180
rect 37714 1708 37854 1718
rect 37714 1596 37854 1606
rect 44620 640 44780 650
rect 44620 470 44780 480
rect 32180 -204 32380 -4
rect 37714 -492 37854 -482
rect 37714 -604 37854 -594
rect 32180 -1044 32380 -844
rect 44620 -1560 44780 -1550
rect 44620 -1730 44780 -1720
rect 40960 -4960 41120 -4950
rect 52620 -4960 52760 2020
rect 58820 2010 58982 2020
rect 41120 -5120 52760 -4960
rect 40960 -5130 41120 -5120
rect 41660 -5380 41820 -5370
rect 41820 -5540 45260 -5380
rect 41660 -5550 41820 -5540
rect 42360 -5720 42520 -5710
rect 42520 -5880 44640 -5720
rect 42360 -5890 42520 -5880
rect 43060 -6140 43220 -6130
rect 43594 -6140 43752 -6139
rect 43220 -6300 44000 -6140
rect 43060 -6310 43220 -6300
rect 34494 -7619 34654 -7609
rect 34654 -7627 36425 -7626
rect 34654 -7629 37771 -7627
rect 34654 -7759 37772 -7629
rect 34494 -7761 37772 -7759
rect 34494 -7763 36425 -7761
rect 34494 -7769 34654 -7763
rect 37602 -8413 37772 -7761
rect 37602 -8529 38085 -8413
rect 34493 -10014 34653 -10010
rect 36514 -10013 37798 -10011
rect 36514 -10014 37845 -10013
rect 34493 -10020 37845 -10014
rect 34653 -10148 37845 -10020
rect 34493 -10170 34653 -10160
rect 37678 -10716 37845 -10148
rect 37676 -10830 38131 -10716
rect 34489 -12417 34649 -12407
rect 36334 -12413 37652 -12412
rect 36334 -12421 37812 -12413
rect 34649 -12555 37812 -12421
rect 34489 -12567 34649 -12557
rect 37616 -12997 37812 -12555
rect 37616 -13118 38090 -12997
rect 34493 -14814 34653 -14804
rect 36314 -14814 37782 -14812
rect 36314 -14824 37784 -14814
rect 34653 -14954 37784 -14824
rect 34493 -14958 37784 -14954
rect 34493 -14964 34653 -14958
rect 37642 -15311 37784 -14958
rect 37642 -15428 38120 -15311
rect 37644 -15436 38120 -15428
rect 34498 -17207 34658 -17197
rect 36414 -17214 37733 -17212
rect 36414 -17220 37734 -17214
rect 34658 -17347 37734 -17220
rect 34498 -17354 37734 -17347
rect 34498 -17357 34658 -17354
rect 36414 -17355 37734 -17354
rect 37518 -17597 37734 -17355
rect 37518 -17720 38100 -17597
rect 34496 -19609 34656 -19599
rect 36334 -19620 37847 -19604
rect 34656 -19749 37847 -19620
rect 34496 -19753 37847 -19749
rect 34496 -19754 37664 -19753
rect 34496 -19759 34656 -19754
rect 37697 -19919 37847 -19753
rect 37697 -20031 38131 -19919
rect 34498 -22011 34658 -22001
rect 36394 -22024 37728 -22018
rect 34658 -22151 37728 -22024
rect 34498 -22158 37728 -22151
rect 34498 -22161 34658 -22158
rect 37554 -22193 37728 -22158
rect 37554 -22317 38113 -22193
rect 34500 -24420 34660 -24410
rect 36354 -24450 38088 -24433
rect 34660 -24560 38088 -24450
rect 34500 -24570 38141 -24560
rect 34572 -24584 38141 -24570
rect 36354 -24590 38141 -24584
rect 43800 -24820 44000 -6300
rect 44460 -15820 44640 -5880
rect 45060 -6820 45260 -5540
rect 58820 -6819 58982 -6809
rect 52900 -6820 58820 -6819
rect 45060 -6980 58820 -6820
rect 58820 -6990 58982 -6980
rect 58820 -15819 58982 -15809
rect 52895 -15820 58820 -15819
rect 44460 -15980 58820 -15820
rect 58820 -15990 58982 -15980
rect 58820 -24819 58982 -24809
rect 43800 -24980 58820 -24820
rect 52899 -24981 58982 -24980
rect 58820 -24990 58982 -24981
<< via2 >>
rect 37714 14806 37854 14908
rect 38200 13360 38360 13520
rect 37714 12606 37854 12708
rect 38880 11180 39040 11320
rect 37714 10406 37854 10508
rect 39580 9020 39740 9180
rect 37714 8206 37854 8308
rect 44620 13680 44780 13840
rect 44620 11480 44780 11640
rect 44620 9280 44780 9440
rect 40280 6920 40440 7080
rect 44620 7080 44780 7240
rect 37714 6006 37854 6108
rect 44620 4880 44780 5040
rect 37714 3806 37854 3908
rect 44620 2680 44780 2840
rect 37714 1606 37854 1708
rect 44620 480 44780 640
rect 37714 -594 37854 -492
rect 44620 -1720 44780 -1560
rect 40960 -5120 41120 -4960
rect 41660 -5540 41820 -5380
rect 42360 -5880 42520 -5720
rect 43060 -6300 43220 -6140
<< metal3 >>
rect 68580 29680 68760 38740
rect 37704 14908 37864 14913
rect 37704 14806 37714 14908
rect 37854 14806 37864 14908
rect 37704 14801 37864 14806
rect 44610 13840 44790 13845
rect 38200 13680 44620 13840
rect 44780 13680 44790 13840
rect 38200 13525 38360 13680
rect 44610 13675 44790 13680
rect 38190 13520 38370 13525
rect 38190 13360 38200 13520
rect 38360 13360 38370 13520
rect 38190 13355 38370 13360
rect 37704 12708 37864 12713
rect 37704 12606 37714 12708
rect 37854 12606 37864 12708
rect 37704 12601 37864 12606
rect 37704 10508 37864 10513
rect 37704 10406 37714 10508
rect 37854 10406 37864 10508
rect 37704 10401 37864 10406
rect 37704 8308 37864 8313
rect 37704 8206 37714 8308
rect 37854 8206 37864 8308
rect 37704 8201 37864 8206
rect 37704 6108 37864 6113
rect 37704 6006 37714 6108
rect 37854 6006 37864 6108
rect 37704 6001 37864 6006
rect 37704 3908 37864 3913
rect 37704 3806 37714 3908
rect 37854 3806 37864 3908
rect 37704 3801 37864 3806
rect 37704 1708 37864 1713
rect 37704 1606 37714 1708
rect 37854 1606 37864 1708
rect 37704 1601 37864 1606
rect 37704 -492 37864 -487
rect 37704 -594 37714 -492
rect 37854 -594 37864 -492
rect 37704 -599 37864 -594
rect 38200 -6740 38360 13355
rect 44610 11640 44790 11645
rect 38880 11480 44620 11640
rect 44780 11480 44790 11640
rect 38880 11475 44790 11480
rect 38880 11460 44700 11475
rect 38880 11345 39040 11460
rect 38870 11320 39050 11345
rect 38870 11180 38880 11320
rect 39040 11180 39050 11320
rect 38870 11175 39050 11180
rect 38450 -6820 38460 -6708
rect 38618 -6820 38628 -6708
rect 38880 -6720 39040 11175
rect 44610 9440 44790 9445
rect 39580 9280 44620 9440
rect 44780 9280 44790 9440
rect 39580 9185 39740 9280
rect 44610 9275 44790 9280
rect 39570 9180 39750 9185
rect 39570 9020 39580 9180
rect 39740 9020 39750 9180
rect 39570 9015 39750 9020
rect 39144 -6820 39154 -6708
rect 39312 -6820 39322 -6708
rect 39580 -6800 39740 9015
rect 44610 7240 44790 7245
rect 40280 7085 44620 7240
rect 40270 7080 44620 7085
rect 44780 7080 44790 7240
rect 40270 6920 40280 7080
rect 40440 6920 40450 7080
rect 44610 7075 44790 7080
rect 40270 6915 40450 6920
rect 39842 -6820 39852 -6708
rect 40010 -6820 40020 -6708
rect 40280 -6800 40440 6915
rect 44610 5040 44790 5045
rect 40960 4880 44620 5040
rect 44780 4880 44790 5040
rect 40960 -4955 41120 4880
rect 44610 4875 44790 4880
rect 44610 2840 44790 2845
rect 41660 2680 44620 2840
rect 44780 2680 44790 2840
rect 40950 -4960 41130 -4955
rect 40950 -5120 40960 -4960
rect 41120 -5120 41130 -4960
rect 40950 -5125 41130 -5120
rect 40536 -6820 40546 -6708
rect 40704 -6820 40714 -6708
rect 40960 -6760 41120 -5125
rect 41660 -5375 41820 2680
rect 44610 2675 44790 2680
rect 44610 640 44790 645
rect 42360 480 44620 640
rect 44780 480 44790 640
rect 41650 -5380 41830 -5375
rect 41650 -5540 41660 -5380
rect 41820 -5540 41830 -5380
rect 41650 -5545 41830 -5540
rect 41226 -6820 41236 -6708
rect 41394 -6820 41404 -6708
rect 41660 -6740 41820 -5545
rect 42360 -5715 42520 480
rect 44610 475 44790 480
rect 44610 -1560 44790 -1555
rect 43060 -1720 44620 -1560
rect 44780 -1720 44790 -1560
rect 42350 -5720 42530 -5715
rect 42350 -5880 42360 -5720
rect 42520 -5880 42530 -5720
rect 42350 -5885 42530 -5880
rect 41920 -6820 41930 -6708
rect 42088 -6820 42098 -6708
rect 42360 -6820 42520 -5885
rect 43060 -6135 43220 -1720
rect 44610 -1725 44790 -1720
rect 43050 -6140 43230 -6135
rect 43050 -6300 43060 -6140
rect 43220 -6300 43230 -6140
rect 43050 -6305 43230 -6300
rect 42618 -6820 42628 -6708
rect 42786 -6820 42796 -6708
rect 43060 -6780 43220 -6305
rect 43312 -6820 43322 -6708
rect 43480 -6820 43490 -6708
<< via3 >>
rect 37714 14806 37854 14908
rect 37714 12606 37854 12708
rect 37714 10406 37854 10508
rect 37714 8206 37854 8308
rect 37714 6006 37854 6108
rect 37714 3806 37854 3908
rect 37714 1606 37854 1708
rect 37714 -594 37854 -492
rect 38460 -6820 38618 -6708
rect 39154 -6820 39312 -6708
rect 39852 -6820 40010 -6708
rect 40546 -6820 40704 -6708
rect 41236 -6820 41394 -6708
rect 41930 -6820 42088 -6708
rect 42628 -6820 42786 -6708
rect 43322 -6820 43480 -6708
<< metal4 >>
rect 37700 14908 43520 14920
rect 37700 14806 37714 14908
rect 37854 14806 43520 14908
rect 37700 14800 43520 14806
rect 37720 12709 42800 12720
rect 37713 12708 42800 12709
rect 37713 12606 37714 12708
rect 37854 12606 42800 12708
rect 37713 12605 42800 12606
rect 37720 12600 42800 12605
rect 37720 10509 42080 10520
rect 37713 10508 42080 10509
rect 37713 10406 37714 10508
rect 37854 10406 42080 10508
rect 37713 10405 42080 10406
rect 37720 10400 42080 10405
rect 37720 8309 41400 8320
rect 37713 8308 41400 8309
rect 37713 8206 37714 8308
rect 37854 8206 41400 8308
rect 37713 8205 41400 8206
rect 37720 8200 41400 8205
rect 37740 6109 40700 6120
rect 37713 6108 40700 6109
rect 37713 6006 37714 6108
rect 37854 6006 40700 6108
rect 37713 6005 40700 6006
rect 37740 6000 40700 6005
rect 37760 3909 40020 3920
rect 37713 3908 40020 3909
rect 37713 3806 37714 3908
rect 37854 3806 40020 3908
rect 37713 3805 40020 3806
rect 37760 3800 40020 3805
rect 37740 1709 39320 1720
rect 37713 1708 39320 1709
rect 37713 1606 37714 1708
rect 37854 1606 39320 1708
rect 37713 1605 39320 1606
rect 37740 1600 39320 1605
rect 37700 -492 38620 -480
rect 37700 -594 37714 -492
rect 37854 -594 38620 -492
rect 37700 -600 38620 -594
rect 38460 -6707 38620 -600
rect 39160 -6707 39320 1600
rect 39860 -6707 40020 3800
rect 38459 -6708 38620 -6707
rect 38459 -6820 38460 -6708
rect 38618 -6780 38620 -6708
rect 39153 -6708 39320 -6707
rect 38618 -6820 38619 -6780
rect 38459 -6821 38619 -6820
rect 39153 -6820 39154 -6708
rect 39312 -6800 39320 -6708
rect 39851 -6708 40020 -6707
rect 39312 -6820 39313 -6800
rect 39153 -6821 39313 -6820
rect 39851 -6820 39852 -6708
rect 40010 -6740 40020 -6708
rect 40540 -6707 40700 6000
rect 41240 -6707 41400 8200
rect 40540 -6708 40705 -6707
rect 40540 -6720 40546 -6708
rect 40010 -6820 40011 -6740
rect 39851 -6821 40011 -6820
rect 40545 -6820 40546 -6720
rect 40704 -6820 40705 -6708
rect 40545 -6821 40705 -6820
rect 41235 -6708 41400 -6707
rect 41235 -6820 41236 -6708
rect 41394 -6720 41400 -6708
rect 41920 -6707 42080 10400
rect 42640 -6707 42800 12600
rect 43340 12540 43520 14800
rect 43340 -6707 43500 12540
rect 41920 -6708 42089 -6707
rect 41920 -6720 41930 -6708
rect 41394 -6820 41395 -6720
rect 41235 -6821 41395 -6820
rect 41929 -6820 41930 -6720
rect 42088 -6820 42089 -6708
rect 41929 -6821 42089 -6820
rect 42627 -6708 42800 -6707
rect 42627 -6820 42628 -6708
rect 42786 -6740 42800 -6708
rect 43321 -6708 43500 -6707
rect 42786 -6820 42787 -6740
rect 42627 -6821 42787 -6820
rect 43321 -6820 43322 -6708
rect 43480 -6740 43500 -6708
rect 43480 -6820 43481 -6740
rect 43321 -6821 43481 -6820
use 8LineSelectOutput04  8LineSelectOutput04_0
timestamp 1700618825
transform 1 0 55900 0 1 0
box 2900 -25000 15779 46870
use 64T64R  x1
timestamp 1700618825
transform 1 0 24980 0 1 -23036
box 13020 -1964 18566 16364
use 8LineSelectInput  x2
timestamp 1700625197
transform -1 0 76136 0 1 -2980
box 27340 400 31536 17916
use 8LineWordInput  x3
timestamp 1700640585
transform 1 0 33036 0 1 -27200
box -2656 1800 1640 22896
use 8LineBitInput  x4
timestamp 1700640585
transform 1 0 -980 0 -1 19196
box 31400 3400 38864 23116
<< labels >>
flabel metal1 48596 2342 48796 2542 0 FreeSans 256 0 0 0 la_data_in96
port 5 nsew
flabel metal1 48595 -2058 48795 -1858 0 FreeSans 256 0 0 0 la_data_in98
flabel metal1 32180 10376 32380 10576 0 FreeSans 256 0 0 0 la_data_in88
port 14 nsew
flabel metal1 32836 -14981 33036 -14781 0 FreeSans 256 0 0 0 la_data_in102
flabel metal1 32835 -17380 33035 -17180 0 FreeSans 256 0 0 0 la_data_in103
port 22 nsew
flabel metal1 32836 -22180 33036 -21980 0 FreeSans 256 0 0 0 la_data_in105
flabel metal1 48160 -1730 48360 -1530 0 FreeSans 256 0 0 0 la_data_in108S
port 30 nsew
flabel metal1 48596 13342 48796 13542 0 FreeSans 256 0 0 0 la_data_in91
port 0 nsew
flabel metal1 48596 11142 48796 11342 0 FreeSans 256 0 0 0 la_data_in92
port 2 nsew
flabel metal1 48596 8942 48796 9142 0 FreeSans 256 0 0 0 la_data_in93
port 3 nsew
flabel metal1 48596 6742 48796 6942 0 FreeSans 256 0 0 0 la_data_in94
port 8 nsew
flabel metal1 48596 4542 48796 4742 0 FreeSans 256 0 0 0 la_data_in95
port 7 nsew
flabel metal1 48576 142 48776 342 0 FreeSans 256 0 0 0 la_data_in97
port 4 nsew
flabel metal1 48596 -2058 48796 -1858 0 FreeSans 256 0 0 0 la_data_in98
port 1 nsew
flabel metal1 32180 14776 32380 14976 0 FreeSans 256 0 0 0 la_data_in90
port 17 nsew
flabel metal1 32180 12576 32380 12776 0 FreeSans 256 0 0 0 la_data_in89
port 16 nsew
flabel metal1 32180 8176 32380 8376 0 FreeSans 256 0 0 0 la_data_in87
port 13 nsew
flabel metal1 32180 5976 32380 6176 0 FreeSans 256 0 0 0 la_data_in86
port 12 nsew
flabel metal1 32180 3776 32380 3976 0 FreeSans 256 0 0 0 la_data_in85
port 11 nsew
flabel metal1 32180 1576 32380 1776 0 FreeSans 256 0 0 0 la_data_in84
port 10 nsew
flabel metal1 32180 -624 32380 -424 0 FreeSans 256 0 0 0 la_data_in83
port 9 nsew
flabel metal1 32836 -7780 33036 -7580 0 FreeSans 256 0 0 0 la_data_in99
port 18 nsew
flabel metal1 32836 -10180 33036 -9980 0 FreeSans 256 0 0 0 la_data_in100
port 19 nsew
flabel metal1 32836 -12580 33036 -12380 0 FreeSans 256 0 0 0 la_data_in101
port 20 nsew
flabel metal1 32836 -14980 33036 -14780 0 FreeSans 256 0 0 0 la_data_in102
port 21 nsew
flabel metal1 32836 -19780 33036 -19580 0 FreeSans 256 0 0 0 la_data_in104
port 23 nsew
flabel metal1 32834 -22180 33034 -21980 0 FreeSans 256 0 0 0 la_data_in105
port 25 nsew
flabel metal1 32836 -24580 33036 -24380 0 FreeSans 256 0 0 0 la_data_in106
port 26 nsew
flabel metal1 30420 -2856 30620 -2656 0 FreeSans 256 0 0 0 la_data_in107B
port 27 nsew
flabel metal2 32180 -1044 32380 -844 0 FreeSans 256 0 0 0 la_data_in108B
port 29 nsew
flabel metal1 30432 -3502 30632 -3302 0 FreeSans 256 0 0 0 v25B
port 31 nsew
flabel metal1 30432 -2388 30632 -2188 0 FreeSans 256 0 0 0 v3B
port 32 nsew
flabel metal2 32180 -204 32380 -4 0 FreeSans 256 0 0 0 v02B
port 33 nsew
flabel metal1 35230 -1694 35430 -1494 0 FreeSans 256 0 0 0 vddB
port 37 nsew
flabel metal1 34080 15572 34280 15772 0 FreeSans 256 0 0 0 vssB
port 38 nsew
flabel metal1 30380 -5568 30580 -5368 0 FreeSans 256 0 0 0 la_data_in107W
port 28 nsew
flabel metal1 30392 -4922 30592 -4722 0 FreeSans 256 0 0 0 v25W
port 34 nsew
flabel metal1 30392 -6034 30592 -5834 0 FreeSans 256 0 0 0 v18W
port 35 nsew
flabel metal1 32940 -25376 33140 -25176 0 FreeSans 256 0 0 0 vssW
port 39 nsew
flabel metal1 32942 -6742 33142 -6542 0 FreeSans 256 0 0 0 vddW
port 40 nsew
flabel metal1 45188 14728 45388 14928 0 FreeSans 256 0 0 0 vdd18SI
port 42 nsew
flabel metal1 46052 14708 46252 14908 0 FreeSans 256 0 0 0 vdd25SI
port 43 nsew
flabel metal1 45186 -2568 45386 -2368 0 FreeSans 256 0 0 0 vssSI
port 44 nsew
flabel metal1 68568 38646 68768 38846 0 FreeSans 256 0 0 0 vssSO
port 46 nsew
flabel metal1 66314 38273 66514 38473 0 FreeSans 256 0 0 0 Gnd
port 47 nsew
flabel metal1 59149 38559 59349 38759 0 FreeSans 256 0 0 0 vssneg
flabel metal1 59150 38559 59350 38759 0 FreeSans 256 0 0 0 vssneg
port 48 nsew
flabel metal1 71478 40048 71678 40248 0 FreeSans 256 0 0 0 la_data_out113
port 49 nsew
flabel metal1 71478 31048 71678 31248 0 FreeSans 256 0 0 0 la_data_out114
port 50 nsew
flabel metal1 71478 22048 71678 22248 0 FreeSans 256 0 0 0 la_data_out115
port 52 nsew
flabel metal1 71478 13048 71678 13248 0 FreeSans 256 0 0 0 la_data_out116
port 53 nsew
flabel metal1 71478 4048 71678 4248 0 FreeSans 256 0 0 0 la_data_out117
port 54 nsew
flabel metal1 71478 -4952 71678 -4752 0 FreeSans 256 0 0 0 la_data_out118
port 55 nsew
flabel metal1 71478 -13952 71678 -13752 0 FreeSans 256 0 0 0 la_data_out119
port 56 nsew
flabel metal1 71478 -22952 71678 -22752 0 FreeSans 256 0 0 0 la_data_out120
port 57 nsew
<< end >>
