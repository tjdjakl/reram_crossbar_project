magic
tech sky130B
magscale 1 2
timestamp 1700694056
<< metal1 >>
rect 13350 696020 13360 696980
rect 14500 696020 14510 696980
rect 26080 696960 28640 696980
rect 26080 696040 26100 696960
rect 28620 696040 28640 696960
rect 68940 696940 71340 697040
rect 13360 682460 14500 696020
rect 26080 695940 28640 696040
rect 68930 696000 68940 696940
rect 71320 696000 71340 696940
rect 68940 695940 71340 696000
rect 120480 696980 122120 697040
rect 120480 696000 120580 696980
rect 122000 696000 122120 696980
rect 120480 695940 122120 696000
rect 26680 693460 28180 695940
rect 69220 695040 71080 695940
rect 120600 694580 121920 695940
rect 118720 693440 118740 693640
rect 118730 693400 118740 693440
rect 119280 693440 120440 693640
rect 122060 693440 122540 693640
rect 123040 693440 123050 693640
rect 119280 693400 119290 693440
rect 28580 693020 41420 693220
rect 41960 693020 41970 693220
rect 71710 692900 71720 692960
rect 71600 692680 71720 692900
rect 72500 692680 72510 692960
rect 17490 692360 17500 692600
rect 18240 692560 18250 692600
rect 18240 692360 26080 692560
rect 28560 692380 36740 692560
rect 37280 692380 37290 692560
rect 28540 691920 38760 692120
rect 39300 691920 39320 692120
rect 26480 685260 28260 691640
rect 68680 691300 69800 691540
rect 68680 691280 69820 691300
rect 68680 691080 68700 691280
rect 69800 691080 69820 691280
rect 120540 685280 122040 692740
rect 26080 685140 28640 685260
rect 120480 685220 122120 685280
rect 26080 684940 26100 685140
rect 26090 684000 26100 684940
rect 28640 684000 28650 685140
rect 120470 683980 120480 685220
rect 122140 683980 122150 685220
rect 12530 681380 12540 681580
rect 12860 681380 13060 681580
rect 14760 681560 15560 681580
rect 14760 681380 15040 681560
rect 15540 681380 15560 681560
rect 13480 680300 14640 680780
rect 13470 679500 13480 680300
rect 14760 679500 14770 680300
rect 441180 666660 442240 671980
rect 556960 666660 557600 668360
rect 441040 666640 442400 666660
rect 441040 666620 442540 666640
rect 441030 664700 441040 666620
rect 442540 664700 442550 666620
rect 556640 666260 557900 666660
rect 556610 664700 556620 666260
rect 557900 664700 557910 666260
rect 4610 646420 4620 646840
rect 4900 646420 4910 646840
rect 5170 645160 5180 645540
rect 5460 645160 5470 645540
rect 4870 644400 4880 644800
rect 5220 644400 5230 644800
rect 579850 641840 579860 642280
rect 580200 641840 580210 642280
rect 580370 640840 580380 641260
rect 580720 640840 580730 641260
rect 580130 640040 580140 640400
rect 580420 640040 580430 640400
rect 54920 273300 55960 273760
rect 36010 272560 36020 273300
rect 37660 272560 55960 273300
rect 7830 222680 7840 223080
rect 8120 222680 8130 223080
rect 7270 219260 7280 219680
rect 7580 219260 7590 219680
rect 6250 217880 6260 218300
rect 6580 217880 6590 218300
rect 7530 217240 7540 217640
rect 7860 217240 7870 217640
rect 5730 216220 5740 216640
rect 6060 216220 6070 216640
rect 6010 215460 6020 215860
rect 6340 215460 6350 215860
rect 194360 103960 240460 104140
rect 240580 103960 240590 104140
rect 194340 91960 244020 92140
rect 244140 91960 244150 92140
rect 50020 87340 51020 88100
rect 36010 86600 36020 87340
rect 37660 86600 51020 87340
rect 490920 83460 527700 83640
rect 527820 83460 527830 83640
rect 194360 79960 247560 80140
rect 247680 79960 247690 80140
rect 490920 74460 531240 74640
rect 531360 74460 531370 74640
rect 194340 67960 251100 68140
rect 251220 67960 251230 68140
rect 158510 65240 158520 66240
rect 159680 66220 159690 66240
rect 159680 65240 159700 66220
rect 490920 65460 534780 65640
rect 534900 65460 534910 65640
rect 158520 62800 159700 65240
rect 158520 62760 187320 62800
rect 158520 61700 186240 62760
rect 187280 61700 187320 62760
rect 158520 61660 187320 61700
rect 158520 58900 159700 61660
rect 454470 61400 454480 61860
rect 455000 61400 455010 61860
rect 454480 59040 455000 61400
rect 150630 58180 150640 58360
rect 150760 58180 156640 58360
rect 444930 58180 444940 58360
rect 445140 58180 451966 58360
rect 490920 56460 538320 56640
rect 538440 56460 538450 56640
rect 147070 55980 147080 56160
rect 147220 55980 156640 56160
rect 194340 55960 254640 56140
rect 254760 55960 254770 56140
rect 441370 55980 441380 56160
rect 441580 55980 451966 56160
rect 173220 54560 173700 54680
rect 173820 54560 173830 54680
rect 468100 54560 468600 54700
rect 468720 54560 468730 54700
rect 50640 53680 52320 53820
rect 143510 53780 143520 53960
rect 143660 53780 156640 53960
rect 437810 53780 437820 53960
rect 438020 53780 451966 53960
rect 50640 53000 50800 53680
rect 52180 53000 52320 53680
rect 50640 51480 52320 53000
rect 173120 52380 174040 52500
rect 174160 52380 174170 52500
rect 468120 52360 468940 52520
rect 469060 52360 469070 52520
rect 139970 51580 139980 51760
rect 140120 51580 156640 51760
rect 434270 51580 434280 51760
rect 434480 51580 451966 51760
rect 173220 50160 174360 50280
rect 174480 50160 174490 50280
rect 468100 50160 469260 50320
rect 469380 50160 469390 50320
rect 50150 49180 50160 49400
rect 50360 49180 50370 49400
rect 136430 49380 136440 49560
rect 136580 49380 156640 49560
rect 430730 49380 430740 49560
rect 430940 49380 451966 49560
rect 52350 47600 52360 48020
rect 53260 47600 53270 48020
rect 173200 47980 174720 48100
rect 174840 47980 174850 48100
rect 468100 47960 469620 48120
rect 469740 47960 469750 48120
rect 490920 47460 541880 47640
rect 542000 47460 542010 47640
rect 132890 47180 132900 47360
rect 133040 47180 156640 47360
rect 427190 47180 427200 47360
rect 427400 47180 451966 47360
rect 173180 45760 175100 45880
rect 175220 45760 175230 45880
rect 468100 45760 470000 45920
rect 470120 45760 470130 45920
rect 129350 44980 129360 45160
rect 129560 44980 156640 45160
rect 423650 44980 423660 45160
rect 423860 44980 451966 45160
rect 194340 43960 258200 44140
rect 258320 43960 258330 44140
rect 173160 43580 175460 43700
rect 175580 43580 175590 43700
rect 468100 43560 470340 43720
rect 470460 43560 470470 43720
rect 125790 42780 125800 42960
rect 126000 42780 156660 42960
rect 420090 42780 420100 42960
rect 420300 42780 451966 42960
rect 173140 41380 176660 41500
rect 176780 41380 176790 41500
rect 468120 41360 473300 41520
rect 473420 41360 473430 41520
rect 152490 40960 152500 41200
rect 152740 41020 155020 41200
rect 447930 41020 447940 41180
rect 448140 41020 449920 41180
rect 152740 40960 152750 41020
rect 169120 40660 170360 40920
rect 158270 40300 158280 40660
rect 158520 40300 170360 40660
rect 464120 40380 465520 40860
rect 452930 39960 452940 40380
rect 453280 39960 465520 40380
rect 154960 39480 157540 39500
rect 449940 39480 452500 39540
rect 154240 39100 157540 39480
rect 445840 39420 452500 39480
rect 445840 39140 445900 39420
rect 446120 39140 452500 39420
rect 445840 39100 452500 39140
rect 28390 38260 28400 38700
rect 28820 38640 28830 38700
rect 154240 38640 154620 39100
rect 154920 39080 157540 39100
rect 449900 39080 452500 39100
rect 155140 39060 157540 39080
rect 155140 39000 157420 39060
rect 28820 38260 154620 38640
rect 490920 38460 545420 38640
rect 545540 38460 545550 38640
rect 154710 35640 154720 35800
rect 154840 35640 157300 35800
rect 449030 35640 449040 35800
rect 449160 35640 452280 35800
rect 155030 33240 155040 33400
rect 155160 33240 157320 33400
rect 449350 33240 449360 33400
rect 449480 33240 452320 33400
rect 194380 31960 261740 32140
rect 261860 31960 261870 32140
rect 155350 30840 155360 31000
rect 155480 30840 157320 31000
rect 449680 30980 452300 31000
rect 449670 30840 449680 30980
rect 449800 30840 452300 30980
rect 490920 29460 548960 29640
rect 549080 29460 549090 29640
rect 155690 28440 155700 28600
rect 155820 28440 157320 28600
rect 450010 28440 450020 28600
rect 450140 28440 452320 28600
rect 156050 26040 156060 26200
rect 156180 26040 157300 26200
rect 450370 26040 450380 26200
rect 450500 26040 452340 26200
rect 156370 23640 156380 23800
rect 156500 23640 157320 23800
rect 450690 23640 450700 23800
rect 450820 23640 452280 23800
rect 156690 21240 156700 21400
rect 156820 21240 157300 21400
rect 451010 21240 451020 21400
rect 451140 21240 452320 21400
rect 50970 20580 50980 21160
rect 52140 20580 52150 21160
rect 50980 19320 52140 20580
rect 490920 20460 552520 20640
rect 552640 20460 552650 20640
rect 194340 19960 265280 20140
rect 265400 19960 265410 20140
rect 52900 18820 72220 19020
rect 72760 18820 72770 19020
rect 156950 18840 156960 19000
rect 157080 18840 157300 19000
rect 451270 18840 451280 19000
rect 451400 18840 452300 19000
rect 48770 18160 48780 18380
rect 49000 18160 50380 18380
rect 162560 18280 163600 18660
rect 457540 18280 458620 18480
rect 158960 18000 163600 18280
rect 453980 18000 458620 18280
rect 80630 17900 80640 17920
rect 52880 17700 80640 17900
rect 81180 17700 81190 17920
rect 51060 16800 52220 17440
rect 51050 16200 51060 16800
rect 52200 16200 52220 16800
rect 51060 16180 52220 16200
<< via1 >>
rect 13360 696020 14500 696980
rect 26100 696040 28620 696960
rect 68940 696000 71320 696940
rect 120580 696000 122000 696980
rect 118740 693400 119280 693640
rect 122540 693440 123040 693640
rect 41420 693020 41960 693220
rect 71720 692680 72500 692960
rect 17500 692360 18240 692600
rect 36740 692380 37280 692560
rect 38760 691920 39300 692120
rect 68700 691080 69800 691280
rect 26100 684000 28640 685140
rect 120480 683980 122140 685220
rect 12540 681380 12860 681580
rect 15040 681380 15540 681560
rect 13480 679500 14760 680300
rect 441040 664700 442540 666620
rect 556620 664700 557900 666260
rect 4620 646420 4900 646840
rect 5180 645160 5460 645540
rect 4880 644400 5220 644800
rect 579860 641840 580200 642280
rect 580380 640840 580720 641260
rect 580140 640040 580420 640400
rect 36020 272560 37660 273300
rect 7840 222680 8120 223080
rect 7280 219260 7580 219680
rect 6260 217880 6580 218300
rect 7540 217240 7860 217640
rect 5740 216220 6060 216640
rect 6020 215460 6340 215860
rect 240460 103960 240580 104140
rect 244020 91960 244140 92140
rect 36020 86600 37660 87340
rect 527700 83460 527820 83640
rect 247560 79960 247680 80140
rect 531240 74460 531360 74640
rect 251100 67960 251220 68140
rect 158520 65240 159680 66240
rect 534780 65460 534900 65640
rect 186240 61700 187280 62760
rect 454480 61400 455000 61860
rect 150640 58180 150760 58360
rect 444940 58180 445140 58360
rect 538320 56460 538440 56640
rect 147080 55980 147220 56160
rect 254640 55960 254760 56140
rect 441380 55980 441580 56160
rect 173700 54560 173820 54680
rect 468600 54560 468720 54700
rect 143520 53780 143660 53960
rect 437820 53780 438020 53960
rect 50800 53000 52180 53680
rect 174040 52380 174160 52500
rect 468940 52360 469060 52520
rect 139980 51580 140120 51760
rect 434280 51580 434480 51760
rect 174360 50160 174480 50280
rect 469260 50160 469380 50320
rect 50160 49180 50360 49400
rect 136440 49380 136580 49560
rect 430740 49380 430940 49560
rect 52360 47600 53260 48020
rect 174720 47980 174840 48100
rect 469620 47960 469740 48120
rect 541880 47460 542000 47640
rect 132900 47180 133040 47360
rect 427200 47180 427400 47360
rect 175100 45760 175220 45880
rect 470000 45760 470120 45920
rect 129360 44980 129560 45160
rect 423660 44980 423860 45160
rect 258200 43960 258320 44140
rect 175460 43580 175580 43700
rect 470340 43560 470460 43720
rect 125800 42780 126000 42960
rect 420100 42780 420300 42960
rect 176660 41380 176780 41500
rect 473300 41360 473420 41520
rect 152500 40960 152740 41200
rect 447940 41020 448140 41180
rect 158280 40300 158520 40660
rect 452940 39960 453280 40380
rect 445900 39140 446120 39420
rect 28400 38260 28820 38700
rect 545420 38460 545540 38640
rect 154720 35640 154840 35800
rect 449040 35640 449160 35800
rect 155040 33240 155160 33400
rect 449360 33240 449480 33400
rect 261740 31960 261860 32140
rect 155360 30840 155480 31000
rect 449680 30840 449800 30980
rect 548960 29460 549080 29640
rect 155700 28440 155820 28600
rect 450020 28440 450140 28600
rect 156060 26040 156180 26200
rect 450380 26040 450500 26200
rect 156380 23640 156500 23800
rect 450700 23640 450820 23800
rect 156700 21240 156820 21400
rect 451020 21240 451140 21400
rect 50980 20580 52140 21160
rect 552520 20460 552640 20640
rect 265280 19960 265400 20140
rect 72220 18820 72760 19020
rect 156960 18840 157080 19000
rect 451280 18840 451400 19000
rect 48780 18160 49000 18380
rect 80640 17700 81180 17920
rect 51060 16200 52200 16800
<< metal2 >>
rect 6420 697060 7720 697070
rect 7720 697040 111560 697060
rect 7720 696980 122040 697040
rect 7720 696020 13360 696980
rect 14500 696960 120580 696980
rect 14500 696040 26100 696960
rect 28620 696940 120580 696960
rect 28620 696040 68940 696940
rect 14500 696020 68940 696040
rect 7720 696000 68940 696020
rect 71320 696000 120580 696940
rect 122000 696000 122040 696980
rect 6420 695990 7720 696000
rect 68940 695990 71320 696000
rect 78240 695980 122040 696000
rect 441340 696340 441580 696350
rect 441340 695890 441580 695900
rect 118740 693640 119280 693650
rect 122540 693640 123040 693650
rect 122540 693430 123040 693440
rect 118740 693390 119280 693400
rect 41420 693220 41960 693230
rect 41420 693010 41960 693020
rect 71720 692960 72500 692970
rect 71720 692670 72500 692680
rect 17500 692600 18240 692610
rect 17500 692350 18240 692360
rect 36740 692560 37280 692580
rect 26100 685140 28640 685150
rect 26100 683990 28640 684000
rect 36740 682920 37280 692380
rect 38760 692120 39300 692130
rect 38760 691910 39300 691920
rect 68700 691280 69800 691290
rect 68700 685140 69800 691080
rect 70080 691180 70300 691190
rect 70080 690950 70300 690960
rect 68700 684030 69800 684040
rect 120480 685220 122140 685230
rect 120480 683970 122140 683980
rect 36740 682050 37280 682060
rect 12540 681580 12860 681590
rect 12540 681370 12860 681380
rect 15040 681560 15540 681570
rect 15040 681370 15540 681380
rect 13480 680300 14760 680310
rect 13480 679490 14760 679500
rect 441380 678960 441580 695890
rect 442140 694380 442380 694390
rect 442140 693930 442380 693940
rect 442140 678940 442340 693930
rect 556960 682100 557160 682110
rect 556960 681670 557160 681680
rect 445980 675980 446520 675990
rect 442420 675800 445980 675980
rect 445980 675730 446520 675740
rect 556960 672720 557140 681670
rect 557640 678480 557840 678490
rect 557640 672720 557840 678060
rect 443680 672320 444220 672330
rect 442420 672120 443680 672320
rect 443680 672030 444220 672040
rect 566960 671140 567500 671150
rect 557860 670940 566960 671140
rect 566960 670930 567500 670940
rect 559840 668820 560380 668830
rect 557880 668640 559840 668820
rect 559840 668630 560380 668640
rect 441040 666620 442540 666630
rect 441040 664690 442540 664700
rect 556620 666260 557900 666270
rect 556620 664690 557900 664700
rect 4620 646840 4900 646850
rect 4620 646410 4900 646420
rect 5180 645540 5460 645550
rect 5180 645150 5460 645160
rect 4880 644800 5220 644810
rect 5220 644400 153760 644800
rect 4880 644390 5220 644400
rect 55760 295660 55960 295670
rect 53940 278680 54240 278690
rect 54240 278500 55260 278680
rect 53940 278490 54240 278500
rect 55060 277960 55260 278500
rect 55760 277980 55960 295280
rect 72220 276400 72760 276410
rect 56020 276200 72220 276400
rect 72220 276190 72760 276200
rect 80640 274100 81180 274110
rect 56020 273900 80640 274100
rect 80640 273890 81180 273900
rect 36020 273300 37660 273310
rect 36020 272550 37660 272560
rect 7840 223080 8120 223090
rect 7840 222670 8120 222680
rect 7280 219680 7580 219690
rect 7280 219250 7580 219260
rect 6260 218300 6580 218310
rect 6260 217870 6580 217880
rect 7540 217640 7860 217650
rect 7860 217240 26360 217640
rect 7540 217230 7860 217240
rect 7560 217220 7840 217230
rect 5740 216640 6060 216650
rect 5740 216210 6060 216220
rect 6020 215860 6340 215870
rect 6340 215460 24260 215860
rect 6020 215450 6340 215460
rect 24000 127290 24260 215460
rect 23900 127280 24440 127290
rect 23900 126690 24440 126700
rect 22720 119840 23260 119850
rect 22720 119250 23260 119260
rect 24000 39280 24260 126690
rect 26100 124710 26360 217240
rect 28560 214050 28820 214060
rect 28400 214040 28820 214050
rect 28780 213520 28820 214040
rect 25980 124700 26520 124710
rect 25980 124110 26520 124120
rect 26100 40200 26360 124110
rect 26100 39910 26360 39920
rect 24000 38990 24260 39000
rect 28400 38700 28820 213520
rect 50980 112340 51180 112350
rect 50240 97100 50440 97110
rect 50240 95000 50440 96900
rect 50980 95040 51180 111960
rect 72220 92080 72760 92090
rect 51200 91880 72220 92080
rect 72220 91870 72760 91880
rect 80640 88400 81180 88410
rect 51160 88200 80640 88400
rect 80640 88190 81180 88200
rect 36020 87340 37660 87350
rect 36020 86590 37660 86600
rect 150640 58360 150760 58370
rect 147080 56160 147220 56170
rect 143520 53960 143660 53970
rect 50800 53680 52180 53690
rect 50800 52990 52180 53000
rect 139980 51760 140120 51770
rect 136440 49560 136580 49570
rect 50160 49400 50360 49410
rect 50160 49170 50360 49180
rect 52360 48020 53260 48030
rect 53260 47600 53280 48000
rect 51640 45120 51880 47580
rect 52360 46760 53280 47600
rect 52360 46200 52400 46760
rect 53220 46200 53280 46760
rect 52360 46140 53280 46200
rect 132900 47360 133040 47370
rect 51640 44910 51880 44920
rect 129360 45160 129560 45170
rect 28400 38250 28820 38260
rect 125800 42960 126000 42970
rect 50980 21160 52140 21170
rect 50980 20570 52140 20580
rect 72220 19020 72760 19030
rect 72220 18810 72760 18820
rect 101080 18400 101620 18410
rect 48780 18380 49000 18390
rect 52880 18180 101080 18380
rect 101620 18180 101640 18380
rect 101080 18170 101620 18180
rect 48780 18150 49000 18160
rect 80640 17920 81180 17930
rect 80640 17690 81180 17700
rect 51060 16800 52200 16810
rect 51060 16190 52200 16200
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125800 400 126000 42780
rect 125816 -800 125928 400
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129360 460 129560 44980
rect 129362 -800 129474 460
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132900 440 133040 47180
rect 132908 -800 133020 440
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136440 420 136580 49380
rect 136454 -800 136566 420
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 139980 440 140120 51580
rect 140000 -800 140112 440
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143520 440 143660 53780
rect 143546 -800 143658 440
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147080 460 147220 55980
rect 150640 480 150760 58180
rect 153360 43420 153760 644400
rect 579860 642280 580200 642290
rect 579860 641830 580200 641840
rect 580380 641260 580720 641270
rect 580380 640830 580720 640840
rect 580140 640400 580420 640410
rect 572100 640380 580140 640400
rect 572100 640040 572140 640380
rect 572680 640040 580140 640380
rect 572140 640030 572680 640040
rect 580140 640030 580420 640040
rect 217320 154380 219140 154390
rect 181080 153300 217320 154280
rect 181080 102740 181520 153300
rect 219140 153320 478160 154280
rect 219140 153300 435500 153320
rect 217320 153270 219140 153280
rect 397780 127220 398040 127240
rect 393780 124620 394080 124630
rect 393780 124110 394080 124120
rect 190820 119820 191240 119830
rect 190820 106160 191240 119280
rect 240460 104140 240580 104150
rect 240460 103880 240580 103960
rect 240460 103860 240581 103880
rect 181080 102460 182060 102740
rect 158520 66240 159680 66250
rect 158520 65230 159680 65240
rect 186240 62760 187280 62770
rect 186240 61690 187280 61700
rect 173700 54680 173820 54690
rect 173700 54550 173820 54560
rect 174040 52500 174160 52510
rect 174040 52370 174160 52380
rect 174360 50280 174480 50290
rect 174360 50150 174480 50160
rect 174720 48100 174840 48110
rect 174720 47970 174840 47980
rect 175100 45880 175220 45890
rect 175100 45750 175220 45760
rect 175460 43700 175580 43710
rect 175460 43570 175580 43580
rect 153360 43160 156660 43420
rect 153320 42380 156720 42540
rect 152500 41200 152740 41210
rect 152500 40950 152740 40960
rect 153320 12940 153440 42380
rect 172800 42200 177100 42340
rect 176660 41500 176780 41510
rect 176660 41370 176780 41380
rect 153880 40700 154000 40710
rect 176980 40680 177100 42200
rect 153880 37980 154000 40560
rect 158280 40660 158520 40670
rect 176980 40550 177100 40560
rect 158280 40290 158520 40300
rect 153880 13480 154000 37840
rect 154720 35800 154840 35810
rect 154720 14300 154840 35640
rect 155040 33400 155160 33410
rect 155040 14920 155160 33240
rect 155360 31000 155480 31010
rect 155360 15500 155480 30840
rect 155700 28600 155820 28610
rect 155700 16040 155820 28440
rect 156060 26200 156180 26210
rect 156060 16500 156180 26040
rect 156380 23800 156500 23810
rect 156380 16960 156500 23640
rect 156700 21400 156820 21410
rect 156700 17380 156820 21240
rect 156960 19000 157080 19010
rect 156960 17780 157080 18840
rect 156960 17640 207500 17780
rect 156700 17240 203940 17380
rect 156380 16820 200400 16960
rect 156060 16360 196860 16500
rect 155700 15900 193300 16040
rect 155360 15360 189760 15500
rect 155040 14780 186220 14920
rect 154720 14160 182660 14300
rect 153880 13330 154000 13340
rect 153320 12790 153440 12800
rect 157720 820 157840 830
rect 154180 740 154300 760
rect 154180 480 154300 600
rect 175460 740 175580 750
rect 171900 720 172020 730
rect 157720 480 157840 680
rect 161260 700 161380 710
rect 161260 480 161380 560
rect 164820 700 164940 710
rect 164820 480 164940 560
rect 168360 700 168480 710
rect 147092 -800 147204 460
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 460 150760 480
rect 150638 -800 150750 460
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157720 460 157842 480
rect 157730 -800 157842 460
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161260 460 161388 480
rect 161276 -800 161388 460
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168360 440 168480 560
rect 171900 480 172020 580
rect 168368 -800 168480 440
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171900 460 172026 480
rect 171914 -800 172026 460
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 440 175580 600
rect 179000 700 179120 710
rect 175460 -800 175572 440
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179000 320 179120 560
rect 182540 480 182660 14160
rect 186100 480 186220 14780
rect 179006 -800 179118 320
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182540 40 182664 480
rect 182552 -800 182664 40
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 20 186220 480
rect 186098 -800 186210 20
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189640 40 189760 15360
rect 193180 480 193300 15900
rect 196740 480 196860 16360
rect 189644 -800 189756 40
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193180 40 193302 480
rect 193190 -800 193302 40
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 160 196860 480
rect 196736 -800 196848 160
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200280 40 200400 16820
rect 200282 -800 200394 40
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203820 240 203940 17240
rect 207380 480 207500 17640
rect 210920 13480 211040 13490
rect 203828 -800 203940 240
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 440 207500 480
rect 207374 -800 207486 440
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 420 211040 13340
rect 214460 12940 214580 12950
rect 210920 -800 211032 420
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214460 20 214580 12800
rect 240461 480 240581 103860
rect 244020 92140 244140 92150
rect 244020 480 244140 91960
rect 247560 80140 247680 80150
rect 214466 -800 214578 20
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240461 415 240582 480
rect 240470 -800 240582 415
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 320 244140 480
rect 244016 -800 244128 320
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247560 420 247680 79960
rect 251100 68140 251220 68150
rect 247562 -800 247674 420
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251100 280 251220 67960
rect 254640 56140 254760 56150
rect 254640 480 254760 55960
rect 258200 44140 258320 44150
rect 251108 -800 251220 280
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254640 320 254766 480
rect 254654 -800 254766 320
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 180 258320 43960
rect 393800 40280 394060 124110
rect 397780 41280 398040 126700
rect 449980 98220 450180 98230
rect 449980 97830 450180 97840
rect 446660 94880 446820 94890
rect 446660 94490 446820 94500
rect 444940 58360 445140 58370
rect 444940 58170 445140 58180
rect 441380 56160 441580 56170
rect 441380 55970 441580 55980
rect 437820 53960 438020 53970
rect 437820 53770 438020 53780
rect 434280 51760 434480 51770
rect 434280 51570 434480 51580
rect 430740 49560 430940 49570
rect 430740 49370 430940 49380
rect 427200 47360 427400 47370
rect 427200 47170 427400 47180
rect 423660 45160 423860 45170
rect 397780 41010 398040 41020
rect 420100 42960 420300 42970
rect 393800 39910 394060 39920
rect 261740 32140 261860 32150
rect 258200 -800 258312 180
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261740 300 261860 31960
rect 265280 20140 265400 20150
rect 265280 480 265400 19960
rect 261746 -800 261858 300
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265280 300 265404 480
rect 265292 -800 265404 300
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420100 400 420300 42780
rect 420134 -800 420246 400
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423660 460 423860 44980
rect 423680 -800 423792 460
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427200 440 427340 47170
rect 430740 480 430880 49370
rect 434280 480 434420 51570
rect 437820 480 437960 53770
rect 441380 480 441520 55970
rect 444940 480 445060 58170
rect 445900 39420 446120 39430
rect 445900 39130 446120 39140
rect 446660 37540 446780 94490
rect 449980 43380 450100 97830
rect 477720 82200 478160 153320
rect 527700 83640 527820 83650
rect 477720 81960 478700 82200
rect 454480 61860 455000 61870
rect 454480 61390 455000 61400
rect 468600 54700 468720 54710
rect 468600 54550 468720 54560
rect 468940 52520 469060 52530
rect 468940 52350 469060 52360
rect 469260 50320 469380 50330
rect 469260 50150 469380 50160
rect 469620 48120 469740 48130
rect 469620 47950 469740 47960
rect 470000 45920 470120 45930
rect 470000 45750 470120 45760
rect 470340 43720 470460 43730
rect 470340 43550 470460 43560
rect 449980 43220 451700 43380
rect 446660 37370 446780 37380
rect 447640 42380 451620 42540
rect 447640 12950 447760 42380
rect 467060 42200 471420 42340
rect 447940 41180 448140 41190
rect 447940 41010 448140 41020
rect 448200 40700 448320 40710
rect 448200 37980 448320 40560
rect 471300 40680 471420 42200
rect 473300 41520 473420 41530
rect 473300 41350 473420 41360
rect 471300 40550 471420 40560
rect 452940 40380 453280 40390
rect 452940 39950 453280 39960
rect 448200 13480 448320 37840
rect 449040 35800 449160 35810
rect 449040 14300 449160 35640
rect 449360 33400 449480 33410
rect 449360 14920 449480 33240
rect 449680 30980 449800 30990
rect 449680 15500 449800 30840
rect 450020 28600 450140 28610
rect 450020 16040 450140 28440
rect 450380 26200 450500 26210
rect 450380 16500 450500 26040
rect 450700 23800 450820 23810
rect 450700 16960 450820 23640
rect 451020 21400 451140 21410
rect 451020 17380 451140 21240
rect 451280 19000 451400 19010
rect 451280 17780 451400 18840
rect 451280 17640 501820 17780
rect 451020 17240 498260 17380
rect 450700 16820 494720 16960
rect 450380 16360 491180 16500
rect 450020 15900 487620 16040
rect 449680 15360 484080 15500
rect 449360 14780 480540 14920
rect 449040 14160 476980 14300
rect 448200 13330 448320 13340
rect 447620 12940 447760 12950
rect 447620 12790 447760 12800
rect 452040 840 452160 850
rect 448500 780 448620 790
rect 427226 -800 427338 440
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430740 420 430884 480
rect 430772 -800 430884 420
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434280 440 434430 480
rect 434318 -800 434430 440
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437820 440 437976 480
rect 437864 -800 437976 440
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441380 460 441522 480
rect 441410 -800 441522 460
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444940 460 445068 480
rect 444956 -800 445068 460
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448500 400 448620 620
rect 470340 800 470460 810
rect 448502 -800 448614 400
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452040 420 452160 680
rect 455580 760 455700 770
rect 455580 480 455700 600
rect 459140 740 459260 750
rect 466220 740 466340 750
rect 452048 -800 452160 420
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455580 360 455706 480
rect 455594 -800 455706 360
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 360 459260 580
rect 462680 720 462800 740
rect 459140 -800 459252 360
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462680 380 462800 560
rect 466220 480 466340 580
rect 469780 640 470340 800
rect 469780 480 469900 640
rect 470340 630 470460 640
rect 473320 800 473440 810
rect 462686 -800 462798 380
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466220 360 466344 480
rect 466232 -800 466344 360
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 380 469900 480
rect 469778 -800 469890 380
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473320 440 473440 640
rect 476860 480 476980 14160
rect 480420 480 480540 14780
rect 473324 -800 473436 440
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476860 40 476982 480
rect 476870 -800 476982 40
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 20 480540 480
rect 480416 -800 480528 20
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483960 40 484080 15360
rect 483962 -800 484074 40
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487500 40 487620 15900
rect 491060 480 491180 16360
rect 487508 -800 487620 40
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 160 491180 480
rect 491054 -800 491166 160
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 40 494720 16820
rect 494600 -800 494712 40
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498140 240 498260 17240
rect 501700 480 501820 17640
rect 505240 13480 505360 13490
rect 505240 480 505360 13340
rect 508780 12940 508900 12950
rect 498146 -800 498258 240
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 440 501820 480
rect 501692 -800 501804 440
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 420 505360 480
rect 505238 -800 505350 420
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508780 20 508900 12800
rect 527700 480 527820 83460
rect 531240 74640 531360 74650
rect 508784 -800 508896 20
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 280 527820 480
rect 527696 -800 527808 280
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531240 400 531360 74460
rect 534780 65640 534900 65650
rect 531242 -800 531354 400
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534780 360 534900 65460
rect 538320 56640 538440 56650
rect 538320 480 538440 56460
rect 541880 47640 542000 47650
rect 534788 -800 534900 360
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538320 320 538446 480
rect 538334 -800 538446 320
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 360 542000 47460
rect 545420 38640 545540 38650
rect 541880 -800 541992 360
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545420 240 545540 38460
rect 548960 29640 549080 29650
rect 548960 480 549080 29460
rect 552520 20640 552640 20650
rect 552520 480 552640 20460
rect 545426 -800 545538 240
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548960 280 549084 480
rect 548972 -800 549084 280
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 300 552640 480
rect 552518 -800 552630 300
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 6420 696000 7720 697060
rect 441340 695900 441580 696340
rect 118740 693400 119280 693640
rect 122540 693440 123040 693640
rect 41420 693020 41960 693220
rect 71720 692680 72500 692960
rect 17500 692360 18240 692600
rect 26100 684000 28640 685140
rect 38760 691920 39300 692120
rect 70080 690960 70300 691180
rect 68700 684040 69800 685140
rect 120480 683980 122140 685220
rect 36740 682060 37280 682920
rect 12540 681380 12860 681580
rect 15040 681380 15540 681560
rect 13480 679500 14760 680300
rect 442140 693940 442380 694380
rect 556960 681680 557160 682100
rect 445980 675740 446520 675980
rect 557640 678060 557840 678480
rect 443680 672040 444220 672320
rect 566960 670940 567500 671140
rect 559840 668640 560380 668820
rect 441040 664700 442540 666620
rect 556620 664700 557900 666260
rect 4620 646420 4900 646840
rect 5180 645160 5460 645540
rect 55760 295280 55960 295660
rect 53940 278500 54240 278680
rect 72220 276200 72760 276400
rect 80640 273900 81180 274100
rect 36020 272560 37660 273300
rect 7840 222680 8120 223080
rect 7280 219260 7580 219680
rect 6260 217880 6580 218300
rect 5740 216220 6060 216640
rect 23900 126700 24440 127280
rect 22720 119260 23260 119840
rect 28400 213520 28780 214040
rect 25980 124120 26520 124700
rect 26100 39920 26360 40200
rect 24000 39000 24260 39280
rect 50980 111960 51180 112340
rect 50240 96900 50440 97100
rect 72220 91880 72760 92080
rect 80640 88200 81180 88400
rect 36020 86600 37660 87340
rect 50800 53000 52180 53680
rect 50160 49180 50360 49400
rect 52400 46200 53220 46760
rect 51640 44920 51880 45120
rect 50980 20580 52140 21160
rect 72220 18820 72760 19020
rect 48780 18160 49000 18380
rect 101080 18180 101620 18400
rect 80640 17700 81180 17920
rect 51060 16200 52200 16800
rect 579860 641840 580200 642280
rect 580380 640840 580720 641260
rect 572140 640040 572680 640380
rect 217320 153280 219140 154380
rect 397780 126700 398040 127220
rect 393780 124120 394080 124620
rect 190820 119280 191240 119820
rect 158520 65240 159680 66240
rect 186240 61700 187280 62760
rect 173700 54560 173820 54680
rect 174040 52380 174160 52500
rect 174360 50160 174480 50280
rect 174720 47980 174840 48100
rect 175100 45760 175220 45880
rect 175460 43580 175580 43700
rect 152500 40960 152740 41200
rect 176660 41380 176780 41500
rect 153880 40560 154000 40700
rect 158280 40300 158520 40660
rect 176980 40560 177100 40680
rect 153880 37840 154000 37980
rect 153880 13340 154000 13480
rect 153320 12800 153440 12940
rect 154180 600 154300 740
rect 157720 680 157840 820
rect 161260 560 161380 700
rect 164820 560 164940 700
rect 168360 560 168480 700
rect 171900 580 172020 720
rect 175460 600 175580 740
rect 179000 560 179120 700
rect 210920 13340 211040 13480
rect 214460 12800 214580 12940
rect 449980 97840 450180 98220
rect 446660 94500 446820 94880
rect 397780 41020 398040 41280
rect 393800 39920 394060 40280
rect 445900 39140 446120 39420
rect 454480 61400 455000 61860
rect 468600 54560 468720 54700
rect 468940 52360 469060 52520
rect 469260 50160 469380 50320
rect 469620 47960 469740 48120
rect 470000 45760 470120 45920
rect 470340 43560 470460 43720
rect 446660 37380 446780 37540
rect 447940 41020 448140 41180
rect 448200 40560 448320 40700
rect 473300 41360 473420 41520
rect 471300 40560 471420 40680
rect 452940 39960 453280 40380
rect 448200 37840 448320 37980
rect 448200 13340 448320 13480
rect 447620 12800 447760 12940
rect 448500 620 448620 780
rect 452040 680 452160 840
rect 455580 600 455700 760
rect 459140 580 459260 740
rect 462680 560 462800 720
rect 466220 580 466340 740
rect 470340 640 470460 800
rect 473320 640 473440 800
rect 505240 13340 505360 13480
rect 508780 12800 508900 12940
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect 6410 697060 7730 697065
rect 6410 696000 6420 697060
rect 7720 696000 7730 697060
rect 6410 695995 7730 696000
rect 17500 692605 18240 702300
rect 41410 693220 41970 693225
rect 41410 693020 41420 693220
rect 41960 693020 41970 693220
rect 41410 693015 41970 693020
rect 71700 692965 72500 702300
rect 122540 693645 123040 702300
rect 414160 696340 415580 702300
rect 441330 696340 441590 696345
rect 414160 695900 441340 696340
rect 441580 695900 441590 696340
rect 441330 695895 441590 695900
rect 442130 694380 442390 694385
rect 467680 694380 469100 702300
rect 442130 693940 442140 694380
rect 442380 693940 469100 694380
rect 442130 693935 442390 693940
rect 118730 693640 119290 693645
rect 118730 693400 118740 693640
rect 119280 693400 119290 693640
rect 122530 693640 123050 693645
rect 122530 693440 122540 693640
rect 123040 693440 123050 693640
rect 122530 693435 123050 693440
rect 118730 693395 119290 693400
rect 71700 692960 72510 692965
rect 71700 692680 71720 692960
rect 72500 692680 72510 692960
rect 71710 692675 72510 692680
rect 17490 692600 18250 692605
rect 17490 692360 17500 692600
rect 18240 692360 18250 692600
rect 17490 692355 18250 692360
rect 38750 692120 39310 692125
rect 38750 691920 38760 692120
rect 39300 691920 39310 692120
rect 38750 691915 39310 691920
rect 70070 691180 70310 691185
rect 70070 690960 70080 691180
rect 70300 690960 70310 691180
rect 70070 690955 70310 690960
rect -800 681580 1700 685242
rect 120470 685220 122150 685225
rect 46800 685200 120480 685220
rect 26080 685140 30900 685200
rect 26080 684000 26100 685140
rect 28640 684000 30900 685140
rect 26080 683960 30900 684000
rect 32900 685140 120480 685200
rect 32900 684040 68700 685140
rect 69800 684040 120480 685140
rect 32900 683980 120480 684040
rect 122140 683980 122150 685220
rect 32900 683960 56100 683980
rect 120470 683975 122150 683980
rect 36730 682920 37290 682925
rect 36730 682060 36740 682920
rect 37280 682060 37290 682920
rect 36730 682055 37290 682060
rect 556950 682100 557170 682105
rect 567640 682100 568900 702300
rect 556950 681680 556960 682100
rect 557160 681680 568900 682100
rect 556950 681675 557170 681680
rect 12530 681580 12870 681585
rect -800 681380 12540 681580
rect 12860 681380 12870 681580
rect -800 680242 1700 681380
rect 12530 681375 12870 681380
rect 15030 681560 15550 681565
rect 15030 681380 15040 681560
rect 15540 681380 15550 681560
rect 441110 681380 441120 681600
rect 441320 681380 441330 681600
rect 15030 681375 15550 681380
rect 13480 680305 30900 680400
rect 13470 680300 30900 680305
rect 13470 679500 13480 680300
rect 14760 679500 30900 680300
rect 13470 679495 30900 679500
rect 13480 679160 30900 679495
rect 32900 679160 32910 680400
rect 441120 678980 441320 681380
rect 441870 679460 441880 679680
rect 442060 679460 442070 679680
rect 441880 678960 442060 679460
rect 582300 678500 584800 682984
rect 557740 678485 584800 678500
rect 557630 678480 584800 678485
rect 557630 678060 557640 678480
rect 557840 678060 584800 678480
rect 557630 678055 557850 678060
rect 582300 677984 584800 678060
rect 445970 675980 446530 675985
rect 445970 675740 445980 675980
rect 446520 675740 446530 675980
rect 445970 675735 446530 675740
rect 556670 674820 556680 675140
rect 556960 674820 556970 675140
rect 556700 672700 556880 674820
rect 557350 673080 557360 673420
rect 557580 673080 557590 673420
rect 557380 672680 557560 673080
rect 443670 672320 444230 672325
rect 443670 672040 443680 672320
rect 444220 672040 444230 672320
rect 443670 672035 444230 672040
rect 566950 671140 567510 671145
rect 566950 670940 566960 671140
rect 567500 670940 567510 671140
rect 566950 670935 567510 670940
rect 559830 668820 560390 668825
rect 559830 668640 559840 668820
rect 560380 668640 560390 668820
rect 559830 668635 560390 668640
rect 442540 666625 510940 666640
rect 441030 666620 510940 666625
rect 441030 664700 441040 666620
rect 442540 664700 510940 666620
rect 512960 666265 557880 666640
rect 512960 666260 557910 666265
rect 512960 664700 556620 666260
rect 557900 664700 557910 666260
rect 441030 664695 442550 664700
rect 556610 664695 557910 664700
rect 41410 660880 41420 661260
rect 41960 660880 70080 661260
rect 70300 660880 118740 661260
rect 119280 660880 445980 661260
rect 446520 660880 566960 661260
rect 567500 660880 567510 661260
rect 38750 658740 38760 659120
rect 39300 658740 443680 659120
rect 444220 658740 559840 659120
rect 560380 658740 560390 659120
rect 436820 656300 436940 656680
rect 437480 656300 543420 656680
rect 543960 656300 543970 656680
rect 433540 652900 433660 653280
rect 434200 652900 535720 653280
rect 536260 652900 536270 653280
rect 2520 651400 3820 651420
rect 2510 650100 2520 651400
rect 3820 650100 3830 651400
rect -800 646860 1660 648642
rect 2520 646860 3820 650100
rect 36730 649560 36740 649940
rect 37280 649920 499600 649940
rect 37280 649560 524120 649920
rect 48680 649540 524120 649560
rect 524660 649540 524670 649920
rect -800 646845 4740 646860
rect -800 646840 4910 646845
rect -800 646420 4620 646840
rect 4900 646420 4910 646840
rect -800 643842 1660 646420
rect 4610 646415 4910 646420
rect 5170 645540 5470 645545
rect 5170 645160 5180 645540
rect 5460 645160 5470 645540
rect 5170 645155 5470 645160
rect 579850 642280 580210 642285
rect 582340 642280 584800 644584
rect 579850 641840 579860 642280
rect 580200 641840 584800 642280
rect 579850 641835 580210 641840
rect 580370 641260 580730 641265
rect 580370 640840 580380 641260
rect 580720 640840 580730 641260
rect 580370 640835 580730 640840
rect 572130 640380 572690 640385
rect 572130 640040 572140 640380
rect 572680 640040 572690 640380
rect 572130 640035 572690 640040
rect 582340 639784 584800 641840
rect -800 637680 1660 638642
rect -800 637460 122800 637680
rect -800 636220 120600 637460
rect 122600 636220 122800 637460
rect -800 636040 122800 636220
rect -800 634280 1660 636040
rect -800 633860 22920 634280
rect 23260 633860 23270 634280
rect -800 633842 7080 633860
rect 1660 633840 7080 633842
rect 582340 631180 584800 634584
rect 577540 631080 584800 631180
rect 577530 629780 577540 631080
rect 578240 629784 584800 631080
rect 578240 629780 583920 629784
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 564240 1660 564242
rect -800 563080 3800 564240
rect 4420 563080 4430 564240
rect -800 561360 1660 563080
rect -800 561280 36020 561360
rect -800 559600 30900 561280
rect 32900 559600 36020 561280
rect -800 559500 36020 559600
rect 37640 559500 37650 560760
rect -800 559442 1660 559500
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 14550 511780 14560 512240
rect 60 511642 14560 511780
rect -800 511530 14560 511642
rect 60 511400 14560 511530
rect 14550 510980 14560 511400
rect 16180 511780 16190 512240
rect 16180 511400 72220 511780
rect 72760 511400 72780 511780
rect 16180 510980 16190 511400
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 60 468420 80640 468540
rect -800 468308 80640 468420
rect 60 468160 80640 468308
rect 81180 468160 81190 468540
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 524110 449580 524120 449960
rect 524660 449830 583760 449960
rect 524660 449718 584800 449830
rect 524660 449580 583760 449718
rect 100 425198 87800 425360
rect -800 425086 87800 425198
rect 100 424980 87800 425086
rect 88340 424980 88350 425360
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 535710 405160 535720 405540
rect 536260 405408 583780 405540
rect 536260 405296 584800 405408
rect 536260 405160 583780 405296
rect 200 381976 94080 382100
rect -800 381864 94080 381976
rect 200 381720 94080 381864
rect 94620 381720 94630 382100
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 543410 358740 543420 359120
rect 543960 358986 583820 359120
rect 543960 358874 584800 358986
rect 543960 358740 583820 358874
rect 60 338754 101080 338900
rect -800 338642 101080 338754
rect 60 338520 101080 338642
rect 101620 338520 101630 338900
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 559830 313520 559840 313900
rect 560380 313764 583720 313900
rect 560380 313652 584800 313764
rect 560380 313520 583720 313652
rect 510950 298360 510960 300300
rect 512980 298360 561320 300300
rect 563340 298360 563350 300300
rect 55750 295660 55970 295665
rect 80 295532 55760 295660
rect -800 295420 55760 295532
rect 80 295280 55760 295420
rect 55960 295280 55970 295660
rect 55750 295275 55970 295280
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 54800 278800 94080 279000
rect 94620 278800 94630 279000
rect 1680 278685 54240 278780
rect 1680 278680 54250 278685
rect 1680 278500 53940 278680
rect 54240 278500 54250 278680
rect 1680 252700 2120 278500
rect 53930 278495 54250 278500
rect 54800 277960 55000 278800
rect 55500 278320 87800 278520
rect 88340 278320 88350 278520
rect 55500 277960 55700 278320
rect 72210 276400 72770 276405
rect 72210 276200 72220 276400
rect 72760 276200 72770 276400
rect 72210 276195 72770 276200
rect 583520 275140 584800 275252
rect 80630 274100 81190 274105
rect 80630 273900 80640 274100
rect 81180 273900 81190 274100
rect 583520 273958 584800 274070
rect 80630 273895 81190 273900
rect 36010 273300 37670 273305
rect 36010 272560 36020 273300
rect 37660 272560 37670 273300
rect 583520 272776 584800 272888
rect 36010 272555 37670 272560
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 566950 269120 566960 269500
rect 567500 269342 583540 269500
rect 567500 269230 584800 269342
rect 567500 269120 583540 269230
rect 60 252510 2120 252700
rect -800 252398 2120 252510
rect 60 252200 2120 252398
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 239360 584800 240030
rect 567530 238640 567540 239360
rect 568100 238640 584800 239360
rect 582340 235230 584800 238640
rect 582340 225230 584800 230030
rect 7830 223080 8130 223085
rect 7830 222680 7840 223080
rect 8120 222680 8130 223080
rect 7830 222675 8130 222680
rect -800 219640 1660 219688
rect 7270 219680 7590 219685
rect 7270 219640 7280 219680
rect -800 219260 7280 219640
rect 7580 219260 7590 219680
rect -800 216640 1660 219260
rect 7270 219255 7590 219260
rect 6250 218300 6590 218305
rect 6250 217880 6260 218300
rect 6580 217880 6590 218300
rect 6250 217875 6590 217880
rect 5730 216640 6070 216645
rect -800 216220 5740 216640
rect 6060 216220 6070 216640
rect -800 214888 1660 216220
rect 3600 214040 4140 216220
rect 5730 216215 6070 216220
rect 28390 214040 28790 214045
rect 3600 213520 28400 214040
rect 28780 213520 28790 214040
rect 28390 213515 28790 213520
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 217310 154380 219150 154385
rect 217310 153280 217320 154380
rect 219140 153280 219150 154380
rect 217310 153275 219150 153280
rect 582340 151460 584800 151630
rect 581070 150020 581080 151460
rect 581640 150020 584800 151460
rect 581080 150000 584800 150020
rect 582340 146830 584800 150000
rect 582340 138500 584800 141630
rect 559400 138440 584800 138500
rect 559400 137200 559480 138440
rect 560320 137200 561320 138440
rect 559400 137080 561320 137200
rect 563340 137080 584800 138440
rect 559400 137040 584800 137080
rect 580912 137038 584800 137040
rect 582340 136830 584800 137038
rect 23890 127280 24450 127285
rect 23890 126700 23900 127280
rect 24440 127240 24450 127280
rect 24440 127225 398020 127240
rect 24440 127220 398050 127225
rect 24440 126700 397780 127220
rect 398040 126700 398050 127220
rect 23890 126695 24450 126700
rect 397770 126695 398050 126700
rect 60 124888 18880 124980
rect -800 124776 18880 124888
rect 60 124640 18880 124776
rect 19420 124640 19430 124980
rect 25970 124700 26530 124705
rect 25970 124120 25980 124700
rect 26520 124660 26540 124700
rect 26520 124620 394120 124660
rect 26520 124120 393780 124620
rect 394080 124120 394120 124620
rect 25970 124115 26530 124120
rect 393770 124115 394090 124120
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect 22710 119840 23270 119845
rect 22710 119260 22720 119840
rect 23260 119820 23270 119840
rect 190810 119820 191250 119825
rect 23260 119280 172280 119820
rect 172620 119280 190820 119820
rect 191240 119280 191260 119820
rect 23260 119260 23270 119280
rect 190810 119275 191250 119280
rect 22710 119255 23270 119260
rect -800 118866 480 118978
rect 50970 112340 51190 112345
rect 18870 111960 18880 112340
rect 19420 111960 50980 112340
rect 51180 111960 51190 112340
rect 50970 111955 51190 111960
rect 454450 105340 454460 105940
rect 455020 105340 559500 105940
rect 560300 105340 560310 105940
rect 567530 103000 567540 103240
rect 445890 102620 445900 102940
rect 446120 102620 567540 103000
rect 568100 102620 568110 103240
rect 449970 98220 450190 98225
rect 572130 98220 572140 98480
rect 449970 97840 449980 98220
rect 450180 97860 572140 98220
rect 572700 98220 572710 98480
rect 572700 97860 572740 98220
rect 450180 97840 572740 97860
rect 449970 97835 450190 97840
rect 50230 97100 50450 97105
rect 560 96900 50240 97100
rect 50440 96900 50450 97100
rect 560 81740 860 96900
rect 50230 96895 50450 96900
rect 49960 96080 94080 96280
rect 94620 96080 94630 96280
rect 49960 95020 50160 96080
rect 50700 95440 87800 95640
rect 88340 95440 88350 95640
rect 50700 95020 50900 95440
rect 583520 95118 584800 95230
rect 446650 94880 446830 94885
rect 446650 94500 446660 94880
rect 446820 94500 464640 94880
rect 465100 94520 577540 94880
rect 578080 94520 578090 94880
rect 465100 94500 578080 94520
rect 446650 94495 446830 94500
rect 72210 92080 72770 92085
rect 72210 91880 72220 92080
rect 72760 91880 72770 92080
rect 72210 91875 72770 91880
rect 80630 88400 81190 88405
rect 80630 88200 80640 88400
rect 81180 88200 81190 88400
rect 80630 88195 81190 88200
rect 36010 87340 37670 87345
rect 36010 86600 36020 87340
rect 37660 86600 37670 87340
rect 36010 86595 37670 86600
rect 488900 85760 489440 94500
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 80 81666 860 81740
rect -800 81554 860 81666
rect 80 81440 860 81554
rect -800 80372 480 80484
rect 482220 80060 482840 81800
rect 454450 79420 454460 80060
rect 455020 79420 488100 80060
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 36010 65220 36020 66360
rect 37660 66240 159700 66360
rect 37660 65240 158520 66240
rect 159680 65240 159700 66240
rect 37660 65220 159700 65240
rect 86420 65200 90860 65220
rect 186220 62760 187320 66220
rect 189180 65020 191640 65240
rect 186220 61700 186240 62760
rect 187280 61700 187320 62760
rect 186220 61660 187320 61700
rect 454470 61860 455010 61865
rect 454470 61400 454480 61860
rect 455000 61400 455010 61860
rect 454470 61395 455010 61400
rect 154180 59740 170700 60020
rect 50790 53680 52190 53685
rect 120590 53680 120600 53820
rect 50790 53000 50800 53680
rect 52180 53000 120600 53680
rect 50790 52995 52190 53000
rect 120590 52960 120600 53000
rect 122560 53680 122570 53820
rect 122560 53000 122600 53680
rect 122560 52960 122570 53000
rect 50150 49400 50370 49405
rect 3880 49180 50160 49400
rect 50360 49180 50370 49400
rect 3880 38480 4280 49180
rect 50150 49175 50370 49180
rect 36010 46140 36020 46800
rect 37640 46760 53280 46800
rect 37640 46200 52400 46760
rect 53220 46200 53280 46760
rect 37640 46140 53280 46200
rect 51630 45120 51890 45125
rect 51630 44920 51640 45120
rect 51880 44920 72220 45120
rect 72760 44920 72770 45120
rect 51630 44915 51890 44920
rect 152490 41200 152750 41205
rect 152490 40960 152500 41200
rect 152740 40960 152750 41200
rect 152490 40955 152750 40960
rect 153870 40700 154010 40705
rect 153870 40560 153880 40700
rect 154000 40560 154010 40700
rect 153870 40555 154010 40560
rect 26090 40200 26370 40205
rect 26090 39920 26100 40200
rect 26360 40080 26370 40200
rect 154180 40080 154400 59740
rect 170500 58120 170700 59740
rect 449400 59740 465920 60020
rect 173040 56760 173540 56920
rect 158270 40660 158530 40665
rect 158270 40300 158280 40660
rect 158520 40300 158530 40660
rect 158270 40295 158530 40300
rect 26360 39920 155000 40080
rect 26090 39915 26370 39920
rect 23990 39280 24270 39285
rect 23990 39000 24000 39280
rect 24260 39180 24270 39280
rect 152490 39180 152500 39260
rect 24260 39020 152500 39180
rect 152740 39020 152750 39260
rect 24260 39000 24270 39020
rect 23990 38995 24270 39000
rect 154180 38660 154400 39920
rect 154180 38500 154940 38660
rect 60 38444 4280 38480
rect -800 38332 4280 38444
rect 60 38260 4280 38332
rect 153870 37980 154010 37985
rect 153870 37840 153880 37980
rect 154000 37840 154010 37980
rect 153870 37835 154010 37840
rect 22910 37380 22920 37740
rect 23240 37540 23260 37740
rect 23240 37380 154940 37540
rect -800 37150 480 37262
rect 158350 37060 158360 37200
rect 158520 37060 158530 37200
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 120570 21240 120580 21260
rect 50940 21160 120580 21240
rect 50940 20580 50980 21160
rect 52140 20580 120580 21160
rect 50940 20560 120580 20580
rect 122580 20560 122590 21260
rect 72210 19020 72770 19025
rect 72210 18820 72220 19020
rect 72760 18820 72770 19020
rect 72210 18815 72770 18820
rect 101070 18400 101630 18405
rect 48770 18380 49010 18385
rect 3740 18160 48780 18380
rect 49000 18160 49010 18380
rect 101070 18180 101080 18400
rect 101620 18180 101630 18400
rect 101070 18175 101630 18180
rect 3740 17060 4060 18160
rect 48770 18155 49010 18160
rect 80630 17920 81190 17925
rect 80630 17700 80640 17920
rect 81180 17700 81190 17920
rect 173420 17900 173540 56760
rect 173700 54685 173820 54700
rect 173690 54680 173830 54685
rect 173690 54560 173700 54680
rect 173820 54560 173830 54680
rect 173690 54555 173830 54560
rect 80630 17695 81190 17700
rect 154180 17780 173540 17900
rect 60 17022 4060 17060
rect -800 16910 4060 17022
rect 60 16840 4060 16910
rect 35990 16160 36000 16860
rect 37620 16840 37630 16860
rect 37620 16800 52240 16840
rect 37620 16200 51060 16800
rect 52200 16200 52240 16800
rect 37620 16160 52240 16200
rect -800 15728 480 15840
rect -800 14546 480 14658
rect 153870 13480 154010 13485
rect -800 13364 480 13476
rect 153870 13340 153880 13480
rect 154000 13340 154010 13480
rect 153870 13335 154010 13340
rect 153310 12940 153450 12945
rect 153310 12800 153320 12940
rect 153440 12800 153450 12940
rect 153310 12795 153450 12800
rect -800 12182 480 12294
rect -800 11000 480 11112
rect -800 9818 480 9930
rect -800 8636 480 8748
rect -800 7454 480 7566
rect -800 6272 480 6384
rect -800 5090 480 5202
rect -800 3908 480 4020
rect -800 2726 480 2838
rect -800 1544 480 1656
rect 154180 745 154300 17780
rect 173700 17640 173820 54555
rect 174040 52505 174160 52520
rect 174030 52500 174170 52505
rect 174030 52380 174040 52500
rect 174160 52380 174170 52500
rect 174030 52375 174170 52380
rect 157720 17520 173820 17640
rect 157720 825 157840 17520
rect 174040 17400 174160 52375
rect 174360 50285 174480 50300
rect 174350 50280 174490 50285
rect 174350 50160 174360 50280
rect 174480 50160 174490 50280
rect 174350 50155 174490 50160
rect 161260 17280 174160 17400
rect 157710 820 157850 825
rect 154170 740 154310 745
rect 154170 600 154180 740
rect 154300 600 154310 740
rect 157710 680 157720 820
rect 157840 680 157850 820
rect 161260 705 161380 17280
rect 174360 17160 174480 50155
rect 174720 48105 174840 48120
rect 174710 48100 174850 48105
rect 174710 47980 174720 48100
rect 174840 47980 174850 48100
rect 174710 47975 174850 47980
rect 164820 17040 174480 17160
rect 164820 705 164940 17040
rect 174720 16900 174840 47975
rect 175100 45885 175220 45900
rect 175090 45880 175230 45885
rect 175090 45760 175100 45880
rect 175220 45760 175230 45880
rect 175090 45755 175230 45760
rect 168360 16780 174840 16900
rect 168360 705 168480 16780
rect 175100 16640 175220 45755
rect 175460 43705 175580 43720
rect 175450 43700 175590 43705
rect 175450 43580 175460 43700
rect 175580 43580 175590 43700
rect 175450 43575 175590 43580
rect 171900 16520 175220 16640
rect 171900 725 172020 16520
rect 175460 745 175580 43575
rect 176650 41500 176790 41505
rect 176650 41380 176660 41500
rect 176780 41380 179120 41500
rect 176650 41375 176790 41380
rect 176970 40680 177110 40685
rect 176970 40560 176980 40680
rect 177100 40560 177110 40680
rect 176970 40555 177110 40560
rect 176980 12940 177100 40555
rect 176970 12800 176980 12940
rect 177100 12800 177110 12940
rect 175450 740 175590 745
rect 171890 720 172030 725
rect 157710 675 157850 680
rect 161250 700 161390 705
rect 154170 595 154310 600
rect 161250 560 161260 700
rect 161380 560 161390 700
rect 161250 555 161390 560
rect 164810 700 164950 705
rect 164810 560 164820 700
rect 164940 560 164950 700
rect 164810 555 164950 560
rect 168350 700 168490 705
rect 168350 560 168360 700
rect 168480 560 168490 700
rect 171890 580 171900 720
rect 172020 580 172030 720
rect 175450 600 175460 740
rect 175580 600 175590 740
rect 179000 705 179120 41380
rect 397770 41280 398050 41285
rect 397770 41020 397780 41280
rect 398040 41180 398050 41280
rect 447930 41180 448150 41185
rect 398040 41020 447940 41180
rect 448140 41020 448150 41180
rect 397770 41015 398050 41020
rect 447930 41015 448150 41020
rect 448190 40700 448330 40705
rect 448190 40560 448200 40700
rect 448320 40560 448330 40700
rect 448190 40555 448330 40560
rect 393790 40280 394070 40285
rect 393790 39920 393800 40280
rect 394060 40080 394070 40280
rect 449400 40080 449620 59740
rect 465720 58300 465920 59740
rect 465660 58120 465920 58300
rect 468060 56760 468440 56920
rect 452930 40380 453290 40385
rect 394060 39920 449960 40080
rect 452930 39960 452940 40380
rect 453280 39960 453290 40380
rect 452930 39955 453290 39960
rect 393790 39915 394070 39920
rect 445890 39420 446130 39425
rect 445890 39140 445900 39420
rect 446120 39140 446130 39420
rect 445890 39135 446130 39140
rect 449400 38660 449620 39920
rect 449400 38500 449900 38660
rect 448190 37980 448330 37985
rect 448190 37840 448200 37980
rect 448320 37840 448330 37980
rect 448190 37835 448330 37840
rect 446650 37540 446790 37545
rect 446650 37380 446660 37540
rect 446780 37380 449900 37540
rect 446650 37375 446790 37380
rect 452910 37060 452920 37200
rect 453280 37080 453290 37200
rect 453280 37060 453340 37080
rect 468320 17900 468440 56760
rect 468590 54700 468730 54705
rect 468590 54560 468600 54700
rect 468720 54560 468730 54700
rect 468590 54555 468730 54560
rect 448500 17780 468440 17900
rect 210910 13480 211050 13485
rect 210910 13340 210920 13480
rect 211040 13340 211050 13480
rect 210910 13335 211050 13340
rect 448190 13480 448330 13485
rect 448190 13340 448200 13480
rect 448320 13340 448330 13480
rect 448190 13335 448330 13340
rect 214450 12940 214590 12945
rect 214450 12800 214460 12940
rect 214580 12800 214590 12940
rect 214450 12795 214590 12800
rect 447610 12940 447770 12945
rect 447610 12800 447620 12940
rect 447760 12800 447770 12940
rect 447610 12795 447770 12800
rect 448500 785 448620 17780
rect 468600 17640 468720 54555
rect 468930 52520 469070 52525
rect 468930 52360 468940 52520
rect 469060 52360 469070 52520
rect 468930 52355 469070 52360
rect 452040 17520 468720 17640
rect 452040 845 452160 17520
rect 468940 17400 469060 52355
rect 583520 50460 584800 50572
rect 469250 50320 469390 50325
rect 469250 50160 469260 50320
rect 469380 50160 469390 50320
rect 469250 50155 469390 50160
rect 455580 17280 469060 17400
rect 452030 840 452170 845
rect 448490 780 448630 785
rect 175450 595 175590 600
rect 178990 700 179130 705
rect 171890 575 172030 580
rect 168350 555 168490 560
rect 178990 560 179000 700
rect 179120 560 179130 700
rect 448490 620 448500 780
rect 448620 620 448630 780
rect 452030 680 452040 840
rect 452160 680 452170 840
rect 455580 765 455700 17280
rect 469260 17160 469380 50155
rect 583520 49278 584800 49390
rect 469610 48120 469750 48125
rect 469610 47960 469620 48120
rect 469740 47960 469750 48120
rect 583520 48096 584800 48208
rect 469610 47955 469750 47960
rect 459140 17040 469380 17160
rect 452030 675 452170 680
rect 455570 760 455710 765
rect 448490 615 448630 620
rect 455570 600 455580 760
rect 455700 600 455710 760
rect 459140 745 459260 17040
rect 469620 16900 469740 47955
rect 583520 46914 584800 47026
rect 469990 45920 470130 45925
rect 469990 45760 470000 45920
rect 470120 45760 470130 45920
rect 469990 45755 470130 45760
rect 462680 16780 469740 16900
rect 455570 595 455710 600
rect 459130 740 459270 745
rect 459130 580 459140 740
rect 459260 580 459270 740
rect 462680 725 462800 16780
rect 470000 16640 470120 45755
rect 470330 43720 470470 43725
rect 470330 43560 470340 43720
rect 470460 43560 470470 43720
rect 470330 43555 470470 43560
rect 466220 16520 470120 16640
rect 466220 745 466340 16520
rect 470340 805 470460 43555
rect 473290 41520 473430 41525
rect 473290 41360 473300 41520
rect 473420 41360 473430 41520
rect 473290 41355 473440 41360
rect 471290 40680 471430 40685
rect 471290 40560 471300 40680
rect 471420 40560 471430 40680
rect 471290 40555 471430 40560
rect 471300 12940 471420 40555
rect 471290 12800 471300 12940
rect 471420 12800 471430 12940
rect 473320 805 473440 41355
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect 583520 16910 584800 17022
rect 583520 15728 584800 15840
rect 583520 14546 584800 14658
rect 505230 13480 505370 13485
rect 505230 13340 505240 13480
rect 505360 13340 505370 13480
rect 583520 13364 584800 13476
rect 505230 13335 505370 13340
rect 508770 12940 508910 12945
rect 508770 12800 508780 12940
rect 508900 12800 508910 12940
rect 508770 12795 508910 12800
rect 583520 12182 584800 12294
rect 583520 11000 584800 11112
rect 583520 9818 584800 9930
rect 583520 8636 584800 8748
rect 583520 7454 584800 7566
rect 583520 6272 584800 6384
rect 583520 5090 584800 5202
rect 583520 3908 584800 4020
rect 583520 2726 584800 2838
rect 583520 1544 584800 1656
rect 470330 800 470470 805
rect 466210 740 466350 745
rect 459130 575 459270 580
rect 462670 720 462810 725
rect 178990 555 179130 560
rect 462670 560 462680 720
rect 462800 560 462810 720
rect 466210 580 466220 740
rect 466340 580 466350 740
rect 470330 640 470340 800
rect 470460 640 470470 800
rect 470330 635 470470 640
rect 473310 800 473450 805
rect 473310 640 473320 800
rect 473440 640 473450 800
rect 473310 635 473450 640
rect 466210 575 466350 580
rect 462670 555 462810 560
rect 179000 540 179120 555
<< via3 >>
rect 6420 696000 7720 697060
rect 41420 693020 41960 693220
rect 118740 693400 119280 693640
rect 38760 691920 39300 692120
rect 70080 690960 70300 691180
rect 30900 683960 32900 685200
rect 36740 682060 37280 682920
rect 15040 681380 15540 681560
rect 441120 681380 441320 681600
rect 30900 679160 32900 680400
rect 441880 679460 442060 679680
rect 445980 675740 446520 675980
rect 556680 674820 556960 675140
rect 557360 673080 557580 673420
rect 443680 672040 444220 672320
rect 566960 670940 567500 671140
rect 559840 668640 560380 668820
rect 510940 664700 512960 666640
rect 41420 660880 41960 661260
rect 70080 660880 70300 661260
rect 118740 660880 119280 661260
rect 445980 660880 446520 661260
rect 566960 660880 567500 661260
rect 38760 658740 39300 659120
rect 443680 658740 444220 659120
rect 559840 658740 560380 659120
rect 436940 656300 437480 656680
rect 543420 656300 543960 656680
rect 433660 652900 434200 653280
rect 535720 652900 536260 653280
rect 2520 650100 3820 651400
rect 36740 649560 37280 649940
rect 524120 649540 524660 649920
rect 5180 645160 5460 645540
rect 580380 640840 580720 641260
rect 572140 640040 572680 640380
rect 120600 636220 122600 637460
rect 22920 633860 23260 634280
rect 577540 629780 578240 631080
rect 3800 563080 4420 564240
rect 30900 559600 32900 561280
rect 36020 559500 37640 560760
rect 14560 510980 16180 512240
rect 72220 511400 72760 511780
rect 80640 468160 81180 468540
rect 524120 449580 524660 449960
rect 87800 424980 88340 425360
rect 535720 405160 536260 405540
rect 94080 381720 94620 382100
rect 543420 358740 543960 359120
rect 101080 338520 101620 338900
rect 559840 313520 560380 313900
rect 510960 298360 512980 300300
rect 561320 298360 563340 300300
rect 94080 278800 94620 279000
rect 87800 278320 88340 278520
rect 72220 276200 72760 276400
rect 80640 273900 81180 274100
rect 36020 272560 37660 273300
rect 566960 269120 567500 269500
rect 567540 238640 568100 239360
rect 7840 222680 8120 223080
rect 6260 217880 6580 218300
rect 217320 153280 219140 154380
rect 581080 150020 581640 151460
rect 559480 137200 560320 138440
rect 561320 137080 563340 138440
rect 18880 124640 19420 124980
rect 172280 119280 172620 119820
rect 18880 111960 19420 112340
rect 454460 105340 455020 105940
rect 559500 105340 560300 105940
rect 445900 102620 446120 102940
rect 567540 102620 568100 103240
rect 572140 97860 572700 98480
rect 94080 96080 94620 96280
rect 87800 95440 88340 95640
rect 464640 94500 465100 94880
rect 577540 94520 578080 94880
rect 72220 91880 72760 92080
rect 80640 88200 81180 88400
rect 36020 86600 37660 87340
rect 454460 79420 455020 80060
rect 36020 65220 37660 66360
rect 454480 61400 455000 61860
rect 120600 52960 122560 53820
rect 36020 46140 37640 46800
rect 72220 44920 72760 45120
rect 152500 40960 152740 41200
rect 153880 40560 154000 40700
rect 158280 40300 158520 40660
rect 152500 39020 152740 39260
rect 153880 37840 154000 37980
rect 22920 37380 23240 37740
rect 158360 37060 158520 37200
rect 120580 20560 122580 21260
rect 72220 18820 72760 19020
rect 101080 18180 101620 18400
rect 80640 17700 81180 17920
rect 36000 16160 37620 16860
rect 153880 13340 154000 13480
rect 153320 12800 153440 12940
rect 176980 12800 177100 12940
rect 448200 40560 448320 40700
rect 452940 39960 453280 40380
rect 445900 39140 446120 39420
rect 448200 37840 448320 37980
rect 452920 37060 453280 37200
rect 210920 13340 211040 13480
rect 448200 13340 448320 13480
rect 214460 12800 214580 12940
rect 447620 12800 447760 12940
rect 471300 12800 471420 12940
rect 505240 13340 505360 13480
rect 508780 12800 508900 12940
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 6419 697060 7721 697061
rect 6419 696000 6420 697060
rect 7720 696000 7721 697060
rect 6419 695999 7721 696000
rect 6420 672940 7720 695999
rect 118739 693640 119281 693641
rect 118739 693400 118740 693640
rect 119280 693400 119281 693640
rect 118739 693399 119281 693400
rect 41419 693220 41961 693221
rect 41419 693020 41420 693220
rect 41960 693020 41961 693220
rect 41419 693019 41961 693020
rect 38759 692120 39301 692121
rect 38759 691920 38760 692120
rect 39300 691920 39301 692120
rect 38759 691919 39301 691920
rect 30899 685200 32901 685201
rect 30899 683960 30900 685200
rect 32900 683960 32901 685200
rect 30899 683959 32901 683960
rect 15039 681560 15541 681561
rect 2520 671760 7720 672940
rect 15020 681380 15040 681560
rect 15540 681380 15560 681560
rect 2520 651401 3820 671760
rect 2519 651400 3821 651401
rect 2519 650100 2520 651400
rect 3820 650100 3821 651400
rect 2519 650099 3821 650100
rect 5179 645540 5461 645541
rect 3980 645160 5180 645540
rect 5460 645160 5461 645540
rect 3980 618720 4440 645160
rect 5179 645159 5461 645160
rect 3980 564241 4420 618720
rect 3799 564240 4421 564241
rect 3799 563080 3800 564240
rect 4420 563080 8200 564240
rect 3799 563079 4421 563080
rect 7760 224000 8200 563080
rect 15020 512241 15560 681380
rect 30900 680401 32900 683959
rect 36739 682920 37281 682921
rect 36739 682060 36740 682920
rect 37280 682060 37281 682920
rect 36739 682059 37281 682060
rect 30899 680400 32901 680401
rect 30899 679160 30900 680400
rect 32900 679160 32901 680400
rect 30899 679159 32901 679160
rect 22919 634280 23261 634281
rect 22919 633860 22920 634280
rect 23260 633860 23261 634280
rect 22720 633859 23261 633860
rect 14559 512240 16181 512241
rect 14559 510980 14560 512240
rect 16180 510980 16181 512240
rect 14559 510979 16181 510980
rect 6220 223200 8200 224000
rect 6220 218300 6660 223200
rect 7760 223080 8200 223200
rect 7760 222680 7840 223080
rect 8120 222680 8200 223080
rect 7839 222679 8121 222680
rect 6220 217880 6260 218300
rect 6580 217880 6660 218300
rect 6259 217879 6581 217880
rect 18879 124980 19421 124981
rect 18879 124640 18880 124980
rect 19420 124640 19421 124980
rect 18879 124639 19421 124640
rect 18880 112341 19420 124639
rect 18879 112340 19421 112341
rect 18879 111960 18880 112340
rect 19420 111960 19421 112340
rect 18879 111959 19421 111960
rect 22720 37740 23260 633859
rect 30900 561281 32900 679159
rect 36740 649941 37280 682059
rect 38760 659121 39300 691919
rect 41420 661261 41960 693019
rect 70079 691180 70301 691181
rect 70079 690960 70080 691180
rect 70300 690960 70301 691180
rect 70079 690959 70301 690960
rect 70080 661261 70300 690959
rect 118740 661261 119280 693399
rect 441119 681600 441321 681601
rect 433660 681380 441120 681600
rect 441320 681380 441321 681600
rect 41419 661260 41961 661261
rect 41419 660880 41420 661260
rect 41960 660880 41961 661260
rect 41419 660879 41961 660880
rect 70079 661260 70301 661261
rect 70079 660880 70080 661260
rect 70300 660880 70301 661260
rect 70079 660879 70301 660880
rect 118739 661260 119281 661261
rect 118739 660880 118740 661260
rect 119280 660880 119281 661260
rect 118739 660879 119281 660880
rect 38759 659120 39301 659121
rect 38759 658740 38760 659120
rect 39300 658740 39301 659120
rect 38759 658739 39301 658740
rect 433660 653281 434200 681380
rect 441119 681379 441321 681380
rect 441879 679680 442061 679681
rect 436940 679460 441880 679680
rect 442060 679460 442080 679680
rect 436940 656681 437480 679460
rect 441879 679459 442061 679460
rect 445979 675980 446521 675981
rect 445979 675740 445980 675980
rect 446520 675740 446521 675980
rect 445979 675739 446521 675740
rect 443679 672320 444221 672321
rect 443679 672040 443680 672320
rect 444220 672040 444221 672320
rect 443679 672039 444221 672040
rect 443680 659121 444220 672039
rect 445980 661261 446520 675739
rect 535720 675140 556980 675160
rect 535720 674820 556680 675140
rect 556960 674820 556980 675140
rect 535720 674800 556980 674820
rect 510939 666640 512961 666641
rect 510939 664700 510940 666640
rect 512960 664700 512961 666640
rect 510939 664699 512961 664700
rect 445979 661260 446521 661261
rect 445979 660880 445980 661260
rect 446520 660880 446521 661260
rect 445979 660879 446521 660880
rect 443679 659120 444221 659121
rect 443679 658740 443680 659120
rect 444220 658740 444221 659120
rect 443679 658739 444221 658740
rect 436939 656680 437481 656681
rect 436939 656300 436940 656680
rect 437480 656300 437481 656680
rect 436939 656299 437481 656300
rect 433659 653280 434201 653281
rect 433659 652900 433660 653280
rect 434200 652900 434201 653280
rect 433659 652899 434201 652900
rect 36739 649940 37281 649941
rect 36739 649560 36740 649940
rect 37280 649560 37281 649940
rect 36739 649559 37281 649560
rect 120599 637460 122601 637461
rect 120599 636220 120600 637460
rect 122600 636220 122601 637460
rect 120599 636219 122601 636220
rect 30899 561280 32901 561281
rect 30899 559600 30900 561280
rect 32900 559600 32901 561280
rect 30899 559599 32901 559600
rect 36019 560760 37641 560761
rect 36019 559500 36020 560760
rect 37640 559500 37660 560760
rect 36019 559499 37660 559500
rect 36020 273301 37660 559499
rect 72219 511780 72761 511781
rect 72219 511400 72220 511780
rect 72760 511400 72761 511780
rect 72219 511399 72761 511400
rect 72220 276401 72760 511399
rect 80639 468540 81181 468541
rect 80639 468160 80640 468540
rect 81180 468160 81181 468540
rect 80639 468159 81181 468160
rect 72219 276400 72761 276401
rect 72219 276200 72220 276400
rect 72760 276200 72761 276400
rect 72219 276199 72761 276200
rect 36019 273300 37661 273301
rect 36019 272560 36020 273300
rect 37660 272560 37661 273300
rect 36019 272559 37661 272560
rect 36020 87341 37660 272559
rect 72220 92081 72760 276199
rect 80640 274101 81180 468159
rect 87799 425360 88341 425361
rect 87799 424980 87800 425360
rect 88340 424980 88341 425360
rect 87799 424979 88341 424980
rect 87800 278521 88340 424979
rect 94079 382100 94621 382101
rect 94079 381720 94080 382100
rect 94620 381720 94621 382100
rect 94079 381719 94621 381720
rect 94080 279001 94620 381719
rect 101079 338900 101621 338901
rect 101079 338520 101080 338900
rect 101620 338520 101621 338900
rect 101079 338519 101621 338520
rect 94079 279000 94621 279001
rect 94079 278800 94080 279000
rect 94620 278800 94621 279000
rect 94079 278799 94621 278800
rect 87799 278520 88341 278521
rect 87799 278320 87800 278520
rect 88340 278320 88341 278520
rect 87799 278319 88341 278320
rect 80639 274100 81181 274101
rect 80639 273900 80640 274100
rect 81180 273900 81181 274100
rect 80639 273899 81181 273900
rect 72219 92080 72761 92081
rect 72219 91880 72220 92080
rect 72760 91880 72761 92080
rect 72219 91879 72761 91880
rect 36019 87340 37661 87341
rect 36019 86600 36020 87340
rect 37660 86600 37661 87340
rect 36019 86599 37661 86600
rect 36020 66361 37660 86599
rect 36019 66360 37661 66361
rect 36019 65220 36020 66360
rect 37660 65220 37661 66360
rect 36019 65219 37661 65220
rect 36020 46801 37660 65219
rect 36019 46800 37660 46801
rect 36019 46140 36020 46800
rect 37640 46140 37660 46800
rect 22720 37380 22920 37740
rect 23240 37380 23260 37740
rect 36000 46139 37641 46140
rect 22919 37379 23241 37380
rect 36000 16861 37640 46139
rect 72220 45121 72760 91879
rect 80640 88401 81180 273899
rect 87800 95641 88340 278319
rect 94080 96281 94620 278799
rect 94079 96280 94621 96281
rect 94079 96080 94080 96280
rect 94620 96080 94621 96280
rect 94079 96079 94621 96080
rect 94080 96000 94620 96079
rect 87799 95640 88341 95641
rect 87799 95440 87800 95640
rect 88340 95440 88341 95640
rect 87799 95439 88341 95440
rect 87800 95420 88340 95439
rect 80639 88400 81181 88401
rect 80639 88200 80640 88400
rect 81180 88200 81181 88400
rect 80639 88199 81181 88200
rect 72219 45120 72761 45121
rect 72219 44920 72220 45120
rect 72760 44920 72761 45120
rect 72219 44919 72761 44920
rect 72220 19021 72760 44919
rect 72219 19020 72761 19021
rect 72219 18820 72220 19020
rect 72760 18820 72761 19020
rect 72219 18819 72761 18820
rect 80640 17921 81180 88199
rect 101080 18401 101620 338519
rect 120600 243960 122600 636219
rect 510940 618760 512940 664699
rect 535720 653281 536260 674800
rect 543420 673420 557600 673440
rect 543420 673080 557360 673420
rect 557580 673080 557600 673420
rect 543420 656681 543960 673080
rect 557359 673079 557581 673080
rect 566959 671140 567501 671141
rect 566959 670940 566960 671140
rect 567500 670940 567501 671140
rect 566959 670939 567501 670940
rect 559839 668820 560381 668821
rect 559839 668640 559840 668820
rect 560380 668640 560381 668820
rect 559839 668639 560381 668640
rect 559840 659121 560380 668639
rect 566960 661261 567500 670939
rect 566959 661260 567501 661261
rect 566959 660880 566960 661260
rect 567500 660880 567501 661260
rect 566959 660879 567501 660880
rect 559839 659120 560381 659121
rect 559839 658740 559840 659120
rect 560380 658740 560381 659120
rect 559839 658739 560381 658740
rect 543419 656680 543961 656681
rect 543419 656300 543420 656680
rect 543960 656300 543961 656680
rect 543419 656299 543961 656300
rect 535719 653280 536261 653281
rect 535719 652900 535720 653280
rect 536260 652900 536261 653280
rect 535719 652899 536261 652900
rect 524119 649920 524661 649921
rect 524119 649540 524120 649920
rect 524660 649540 524661 649920
rect 524119 649539 524661 649540
rect 510940 547060 512980 618760
rect 510960 300301 512980 547060
rect 524120 449961 524660 649539
rect 524119 449960 524661 449961
rect 524119 449580 524120 449960
rect 524660 449580 524661 449960
rect 524119 449579 524661 449580
rect 535720 405541 536260 652899
rect 535719 405540 536261 405541
rect 535719 405160 535720 405540
rect 536260 405160 536261 405540
rect 535719 405159 536261 405160
rect 543420 359121 543960 656299
rect 543419 359120 543961 359121
rect 543419 358740 543420 359120
rect 543960 358740 543961 359120
rect 543419 358739 543961 358740
rect 559840 313901 560380 658739
rect 559839 313900 560381 313901
rect 559839 313520 559840 313900
rect 560380 313520 560381 313900
rect 559839 313519 560381 313520
rect 510959 300300 512981 300301
rect 510959 298360 510960 300300
rect 512980 298360 512981 300300
rect 510959 298359 512981 298360
rect 561319 300300 563341 300301
rect 561319 298360 561320 300300
rect 563340 298360 563341 300300
rect 561319 298359 563341 298360
rect 120580 107500 122600 243960
rect 217319 154380 219141 154381
rect 217319 153280 217320 154380
rect 219140 153280 219141 154380
rect 217319 153279 219141 153280
rect 561320 138441 563340 298359
rect 566960 269501 567500 660879
rect 580379 641260 580721 641261
rect 580379 640840 580380 641260
rect 580720 640840 581420 641260
rect 580379 640839 580721 640840
rect 572139 640380 572681 640381
rect 572139 640040 572140 640380
rect 572680 640040 572681 640380
rect 572139 639959 572681 640040
rect 566959 269500 567501 269501
rect 566959 269120 566960 269500
rect 567500 269120 567501 269500
rect 566959 269119 567501 269120
rect 567539 239360 568101 239361
rect 567539 238640 567540 239360
rect 568100 238640 568101 239360
rect 567539 238639 568101 238640
rect 559479 138440 560321 138441
rect 559479 137200 559480 138440
rect 560320 137200 560321 138440
rect 559479 137199 560321 137200
rect 561319 138440 563341 138441
rect 172279 119820 172621 119821
rect 172220 119280 172280 119820
rect 172620 119280 172621 119820
rect 172220 119279 172621 119280
rect 120580 53820 122580 107500
rect 172220 58120 172620 119279
rect 454459 105940 455021 105941
rect 454459 105340 454460 105940
rect 455020 105340 455021 105940
rect 454459 105339 455021 105340
rect 559480 105940 560320 137199
rect 561319 137080 561320 138440
rect 563340 137080 563341 138440
rect 561319 137079 563341 137080
rect 559480 105340 559500 105940
rect 560300 105340 560320 105940
rect 445900 102941 446120 103000
rect 445899 102940 446121 102941
rect 445899 102620 445900 102940
rect 446120 102620 446121 102940
rect 445899 102619 446121 102620
rect 120580 52960 120600 53820
rect 122560 52960 122580 53820
rect 120580 21261 122580 52960
rect 158360 41540 158640 41560
rect 158280 41380 158640 41540
rect 152499 41200 152741 41201
rect 152499 40960 152500 41200
rect 152740 40960 152741 41200
rect 152499 40959 152741 40960
rect 152500 39261 152740 40959
rect 153879 40700 154001 40701
rect 153879 40560 153880 40700
rect 154000 40560 154980 40700
rect 158280 40661 158520 41380
rect 158279 40660 158521 40661
rect 153879 40559 154001 40560
rect 158279 40300 158280 40660
rect 158520 40300 158521 40660
rect 158279 40299 158521 40300
rect 152499 39260 152741 39261
rect 152499 39020 152500 39260
rect 152740 39020 152741 39260
rect 152499 39019 152741 39020
rect 153879 37980 154001 37981
rect 153879 37840 153880 37980
rect 154000 37840 154900 37980
rect 153879 37839 154001 37840
rect 158280 37201 158520 40299
rect 445900 39421 446120 102619
rect 454460 80061 455020 105339
rect 559480 105320 560320 105340
rect 567540 103241 568100 238639
rect 572140 105200 572680 639959
rect 577539 631080 578241 631081
rect 577539 629780 577540 631080
rect 578240 629780 578241 631080
rect 577539 629779 578241 629780
rect 567539 103240 568101 103241
rect 567539 102620 567540 103240
rect 568100 102620 568101 103240
rect 567539 102619 568101 102620
rect 572140 98481 572700 105200
rect 572139 98480 572701 98481
rect 572139 97860 572140 98480
rect 572700 97860 572701 98480
rect 572139 97859 572701 97860
rect 464660 94881 465060 94900
rect 577540 94881 578080 629779
rect 581080 151461 581420 640840
rect 581079 151460 581641 151461
rect 581079 150020 581080 151460
rect 581640 150020 581641 151460
rect 581079 150019 581641 150020
rect 464639 94880 465101 94881
rect 464639 94500 464640 94880
rect 465100 94500 465101 94880
rect 577539 94880 578081 94881
rect 577539 94520 577540 94880
rect 578080 94520 578081 94880
rect 577539 94519 578081 94520
rect 464639 94499 465101 94500
rect 454459 80060 455021 80061
rect 454459 79420 454460 80060
rect 455020 79420 455021 80060
rect 454459 79419 455021 79420
rect 454460 61860 455020 79419
rect 454460 61400 454480 61860
rect 455000 61400 455020 61860
rect 454460 61380 455020 61400
rect 464660 58140 465060 94499
rect 448199 40700 448321 40701
rect 448199 40560 448200 40700
rect 448320 40560 449960 40700
rect 448199 40559 448321 40560
rect 452920 40380 453300 41560
rect 452920 39960 452940 40380
rect 453280 39960 453300 40380
rect 445899 39420 446121 39421
rect 445899 39140 445900 39420
rect 446120 39140 446121 39420
rect 445899 39139 446121 39140
rect 448199 37980 448321 37981
rect 448199 37840 448200 37980
rect 448320 37840 449900 37980
rect 448199 37839 448321 37840
rect 452920 37201 453300 39960
rect 158280 37200 158521 37201
rect 158280 37060 158360 37200
rect 158520 37060 158521 37200
rect 158359 37059 158521 37060
rect 452919 37200 453300 37201
rect 452919 37060 452920 37200
rect 453280 37060 453300 37200
rect 452919 37059 453281 37060
rect 120579 21260 122581 21261
rect 120579 20560 120580 21260
rect 122580 20560 122581 21260
rect 120579 20559 122581 20560
rect 101079 18400 101621 18401
rect 101079 18180 101080 18400
rect 101620 18180 101621 18400
rect 101079 18179 101621 18180
rect 80639 17920 81181 17921
rect 80639 17700 80640 17920
rect 81180 17700 81181 17920
rect 80639 17699 81181 17700
rect 35999 16860 37640 16861
rect 35999 16160 36000 16860
rect 37620 16160 37640 16860
rect 35999 16159 37621 16160
rect 120580 10140 122580 20559
rect 153879 13480 154001 13481
rect 210919 13480 211041 13481
rect 153879 13340 153880 13480
rect 154000 13340 210920 13480
rect 211040 13340 211041 13480
rect 153879 13339 154001 13340
rect 210919 13339 211041 13340
rect 448199 13480 448321 13481
rect 505239 13480 505361 13481
rect 448199 13340 448200 13480
rect 448320 13340 505240 13480
rect 505360 13340 505361 13480
rect 448199 13339 448321 13340
rect 505239 13339 505361 13340
rect 153319 12940 153441 12941
rect 176979 12940 177101 12941
rect 214459 12940 214581 12941
rect 153319 12800 153320 12940
rect 153440 12800 176980 12940
rect 177100 12800 214460 12940
rect 214580 12800 214581 12940
rect 153319 12799 153441 12800
rect 176979 12799 177101 12800
rect 214459 12799 214581 12800
rect 447619 12940 447761 12941
rect 471299 12940 471421 12941
rect 508779 12940 508901 12941
rect 447619 12800 447620 12940
rect 447760 12800 471300 12940
rect 471420 12800 508780 12940
rect 508900 12800 508901 12940
rect 447619 12799 447761 12800
rect 471299 12799 471421 12800
rect 508779 12799 508901 12800
<< via4 >>
rect 217320 153280 219140 154380
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 217320 154404 219140 702300
rect 217296 154380 219164 154404
rect 217296 153280 217320 154380
rect 219140 153280 219164 154380
rect 217296 153256 219164 153280
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use 2-1MUX  2-1MUX_0 ~/ReRAM_Crossbar_Project/magic
timestamp 1700640585
transform -1 0 27804 0 1 690920
box -936 600 1824 2716
use 2-1MUX  2-1MUX_1
timestamp 1700640585
transform -1 0 52144 0 1 16720
box -936 600 1824 2716
use 02Compute  02Compute_0 ~/ReRAM_Crossbar_Project/magic
timestamp 1700640585
transform 1 0 124446 0 1 43400
box 30380 -25400 70090 70482
use 04Compute  04Compute_0 ~/ReRAM_Crossbar_Project/magic
timestamp 1700640585
transform 1 0 419426 0 1 43400
box 30380 -25400 71679 46870
use 4T4R  4T4R_0 ~/ReRAM_Crossbar_Project/magic
timestamp 1700618825
transform -1 0 558480 0 1 667406
box 462 854 1840 5424
use 4T4R  4T4R_1
timestamp 1700618825
transform -1 0 56600 0 1 272666
box 462 854 1840 5424
use 4T4RLarge  4T4RLarge_0 ~/ReRAM_Crossbar_Project/magic
timestamp 1700640568
transform -1 0 447014 0 1 672750
box 4508 -970 5974 6336
use 4T4RLarge  4T4RLarge_1
timestamp 1700640568
transform -1 0 55854 0 1 88830
box 4508 -970 5974 6336
use Buffer  Buffer_0 ~/ReRAM_Crossbar_Project/magic
timestamp 1700618825
transform 1 0 118522 0 1 691260
box 1858 1360 3698 3442
use Buffer  Buffer_1
timestamp 1700618825
transform -1 0 16718 0 1 679200
box 1858 1360 3698 3442
use oneBitADC  oneBitADC_0 ~/ReRAM_Crossbar_Project/magic
timestamp 1700618825
transform 1 0 67504 0 1 690452
box 656 288 4296 4810
use oneBitADC  oneBitADC_1
timestamp 1700618825
transform -1 0 54456 0 1 46952
box 656 288 4296 4810
use vDivider_02  vDivider_02_0 ~/ReRAM_Crossbar_Project/magic
timestamp 1697725649
transform 1 0 4573 0 1 643674
box -53 546 1014 3339
use vDivider_3  vDivider_3_0 ~/ReRAM_Crossbar_Project/magic
timestamp 1697725649
transform 1 0 5746 0 1 214786
box -106 494 958 3686
use vDivider_04  vDivider_04_0 ~/ReRAM_Crossbar_Project/magic
timestamp 1697725317
transform 1 0 579813 0 1 639294
box -53 546 1006 3139
use vDivider_25  vDivider_25_0 ~/ReRAM_Crossbar_Project/magic
timestamp 1700613895
transform 1 0 7286 0 1 216568
box -106 492 958 6686
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
