magic
tech sky130B
magscale 1 2
timestamp 1688980957
use sky130_fd_pr__dfl1sd__example_55959141808190  sky130_fd_pr__dfl1sd__example_55959141808190_0
timestamp 1688980957
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808190  sky130_fd_pr__dfl1sd__example_55959141808190_1
timestamp 1688980957
transform 1 0 50 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 3514182
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3513260
<< end >>
