magic
tech sky130B
magscale 1 2
timestamp 1700618825
<< pwell >>
rect -1765 -3733 1765 3733
<< psubdiff >>
rect -1729 3663 -1633 3697
rect 1633 3663 1729 3697
rect -1729 3601 -1695 3663
rect 1695 3601 1729 3663
rect -1729 -3663 -1695 -3601
rect 1695 -3663 1729 -3601
rect -1729 -3697 -1633 -3663
rect 1633 -3697 1729 -3663
<< psubdiffcont >>
rect -1633 3663 1633 3697
rect -1729 -3601 -1695 3601
rect 1695 -3601 1729 3601
rect -1633 -3697 1633 -3663
<< poly >>
rect -1599 -3517 -1533 -3137
rect -1599 -3551 -1583 -3517
rect -1549 -3551 -1533 -3517
rect -1599 -3567 -1533 -3551
rect 1533 -3517 1599 -3137
rect 1533 -3551 1549 -3517
rect 1583 -3551 1599 -3517
rect 1533 -3567 1599 -3551
<< polycont >>
rect -1583 -3551 -1549 -3517
rect 1549 -3551 1583 -3517
<< npolyres >>
rect -1599 3501 -1425 3567
rect -1599 -3137 -1533 3501
rect -1491 -2967 -1425 3501
rect -1383 3501 -1209 3567
rect -1383 -2967 -1317 3501
rect -1491 -3033 -1317 -2967
rect -1275 -2967 -1209 3501
rect -1167 3501 -993 3567
rect -1167 -2967 -1101 3501
rect -1275 -3033 -1101 -2967
rect -1059 -2967 -993 3501
rect -951 3501 -777 3567
rect -951 -2967 -885 3501
rect -1059 -3033 -885 -2967
rect -843 -2967 -777 3501
rect -735 3501 -561 3567
rect -735 -2967 -669 3501
rect -843 -3033 -669 -2967
rect -627 -2967 -561 3501
rect -519 3501 -345 3567
rect -519 -2967 -453 3501
rect -627 -3033 -453 -2967
rect -411 -2967 -345 3501
rect -303 3501 -129 3567
rect -303 -2967 -237 3501
rect -411 -3033 -237 -2967
rect -195 -2967 -129 3501
rect -87 3501 87 3567
rect -87 -2967 -21 3501
rect -195 -3033 -21 -2967
rect 21 -2967 87 3501
rect 129 3501 303 3567
rect 129 -2967 195 3501
rect 21 -3033 195 -2967
rect 237 -2967 303 3501
rect 345 3501 519 3567
rect 345 -2967 411 3501
rect 237 -3033 411 -2967
rect 453 -2967 519 3501
rect 561 3501 735 3567
rect 561 -2967 627 3501
rect 453 -3033 627 -2967
rect 669 -2967 735 3501
rect 777 3501 951 3567
rect 777 -2967 843 3501
rect 669 -3033 843 -2967
rect 885 -2967 951 3501
rect 993 3501 1167 3567
rect 993 -2967 1059 3501
rect 885 -3033 1059 -2967
rect 1101 -2967 1167 3501
rect 1209 3501 1383 3567
rect 1209 -2967 1275 3501
rect 1101 -3033 1275 -2967
rect 1317 -2967 1383 3501
rect 1425 3501 1599 3567
rect 1425 -2967 1491 3501
rect 1317 -3033 1491 -2967
rect 1533 -3137 1599 3501
<< locali >>
rect -1729 3663 -1633 3697
rect 1633 3663 1729 3697
rect -1729 3601 -1695 3663
rect 1695 3601 1729 3663
rect -1599 -3551 -1583 -3517
rect -1549 -3551 -1533 -3517
rect 1533 -3551 1549 -3517
rect 1583 -3551 1599 -3517
rect -1729 -3663 -1695 -3601
rect 1695 -3663 1729 -3601
rect -1729 -3697 -1633 -3663
rect 1633 -3697 1729 -3663
<< properties >>
string FIXED_BBOX -1712 -3680 1712 3680
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.330 l 33 m 1 nx 30 wmin 0.330 lmin 1.650 rho 48.2 val 147.692k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 1 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
