magic
tech sky130B
magscale 1 2
timestamp 1700538807
<< pwell >>
rect -1333 -2203 1333 2203
<< psubdiff >>
rect -1297 2133 -1201 2167
rect 1201 2133 1297 2167
rect -1297 2071 -1263 2133
rect 1263 2071 1297 2133
rect -1297 -2133 -1263 -2071
rect 1263 -2133 1297 -2071
rect -1297 -2167 -1201 -2133
rect 1201 -2167 1297 -2133
<< psubdiffcont >>
rect -1201 2133 1201 2167
rect -1297 -2071 -1263 2071
rect 1263 -2071 1297 2071
rect -1201 -2167 1201 -2133
<< poly >>
rect -1167 -1987 -1101 -1607
rect -1167 -2021 -1151 -1987
rect -1117 -2021 -1101 -1987
rect -1167 -2037 -1101 -2021
rect 1101 -1987 1167 -1607
rect 1101 -2021 1117 -1987
rect 1151 -2021 1167 -1987
rect 1101 -2037 1167 -2021
<< polycont >>
rect -1151 -2021 -1117 -1987
rect 1117 -2021 1151 -1987
<< npolyres >>
rect -1167 1971 -993 2037
rect -1167 -1607 -1101 1971
rect -1059 -1437 -993 1971
rect -951 1971 -777 2037
rect -951 -1437 -885 1971
rect -1059 -1503 -885 -1437
rect -843 -1437 -777 1971
rect -735 1971 -561 2037
rect -735 -1437 -669 1971
rect -843 -1503 -669 -1437
rect -627 -1437 -561 1971
rect -519 1971 -345 2037
rect -519 -1437 -453 1971
rect -627 -1503 -453 -1437
rect -411 -1437 -345 1971
rect -303 1971 -129 2037
rect -303 -1437 -237 1971
rect -411 -1503 -237 -1437
rect -195 -1437 -129 1971
rect -87 1971 87 2037
rect -87 -1437 -21 1971
rect -195 -1503 -21 -1437
rect 21 -1437 87 1971
rect 129 1971 303 2037
rect 129 -1437 195 1971
rect 21 -1503 195 -1437
rect 237 -1437 303 1971
rect 345 1971 519 2037
rect 345 -1437 411 1971
rect 237 -1503 411 -1437
rect 453 -1437 519 1971
rect 561 1971 735 2037
rect 561 -1437 627 1971
rect 453 -1503 627 -1437
rect 669 -1437 735 1971
rect 777 1971 951 2037
rect 777 -1437 843 1971
rect 669 -1503 843 -1437
rect 885 -1437 951 1971
rect 993 1971 1167 2037
rect 993 -1437 1059 1971
rect 885 -1503 1059 -1437
rect 1101 -1607 1167 1971
<< locali >>
rect -1297 2133 -1201 2167
rect 1201 2133 1297 2167
rect -1297 2071 -1263 2133
rect 1263 2071 1297 2133
rect -1167 -2021 -1151 -1987
rect -1117 -2021 -1101 -1987
rect 1101 -2021 1117 -1987
rect 1151 -2021 1167 -1987
rect -1297 -2133 -1263 -2071
rect 1263 -2133 1297 -2071
rect -1297 -2167 -1201 -2133
rect 1201 -2167 1297 -2133
<< properties >>
string FIXED_BBOX -1280 -2150 1280 2150
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.33 l 17.7 m 1 nx 22 wmin 0.330 lmin 1.650 rho 48.2 val 59.115k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 1 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
