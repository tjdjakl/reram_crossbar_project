magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect 0 0 294 1072
<< pmos >>
rect 89 36 119 1036
rect 175 36 205 1036
<< pdiff >>
rect 36 985 89 1036
rect 36 951 44 985
rect 78 951 89 985
rect 36 913 89 951
rect 36 879 44 913
rect 78 879 89 913
rect 36 841 89 879
rect 36 807 44 841
rect 78 807 89 841
rect 36 769 89 807
rect 36 735 44 769
rect 78 735 89 769
rect 36 697 89 735
rect 36 663 44 697
rect 78 663 89 697
rect 36 625 89 663
rect 36 591 44 625
rect 78 591 89 625
rect 36 553 89 591
rect 36 519 44 553
rect 78 519 89 553
rect 36 481 89 519
rect 36 447 44 481
rect 78 447 89 481
rect 36 409 89 447
rect 36 375 44 409
rect 78 375 89 409
rect 36 337 89 375
rect 36 303 44 337
rect 78 303 89 337
rect 36 265 89 303
rect 36 231 44 265
rect 78 231 89 265
rect 36 193 89 231
rect 36 159 44 193
rect 78 159 89 193
rect 36 121 89 159
rect 36 87 44 121
rect 78 87 89 121
rect 36 36 89 87
rect 119 985 175 1036
rect 119 951 130 985
rect 164 951 175 985
rect 119 913 175 951
rect 119 879 130 913
rect 164 879 175 913
rect 119 841 175 879
rect 119 807 130 841
rect 164 807 175 841
rect 119 769 175 807
rect 119 735 130 769
rect 164 735 175 769
rect 119 697 175 735
rect 119 663 130 697
rect 164 663 175 697
rect 119 625 175 663
rect 119 591 130 625
rect 164 591 175 625
rect 119 553 175 591
rect 119 519 130 553
rect 164 519 175 553
rect 119 481 175 519
rect 119 447 130 481
rect 164 447 175 481
rect 119 409 175 447
rect 119 375 130 409
rect 164 375 175 409
rect 119 337 175 375
rect 119 303 130 337
rect 164 303 175 337
rect 119 265 175 303
rect 119 231 130 265
rect 164 231 175 265
rect 119 193 175 231
rect 119 159 130 193
rect 164 159 175 193
rect 119 121 175 159
rect 119 87 130 121
rect 164 87 175 121
rect 119 36 175 87
rect 205 985 258 1036
rect 205 951 216 985
rect 250 951 258 985
rect 205 913 258 951
rect 205 879 216 913
rect 250 879 258 913
rect 205 841 258 879
rect 205 807 216 841
rect 250 807 258 841
rect 205 769 258 807
rect 205 735 216 769
rect 250 735 258 769
rect 205 697 258 735
rect 205 663 216 697
rect 250 663 258 697
rect 205 625 258 663
rect 205 591 216 625
rect 250 591 258 625
rect 205 553 258 591
rect 205 519 216 553
rect 250 519 258 553
rect 205 481 258 519
rect 205 447 216 481
rect 250 447 258 481
rect 205 409 258 447
rect 205 375 216 409
rect 250 375 258 409
rect 205 337 258 375
rect 205 303 216 337
rect 250 303 258 337
rect 205 265 258 303
rect 205 231 216 265
rect 250 231 258 265
rect 205 193 258 231
rect 205 159 216 193
rect 250 159 258 193
rect 205 121 258 159
rect 205 87 216 121
rect 250 87 258 121
rect 205 36 258 87
<< pdiffc >>
rect 44 951 78 985
rect 44 879 78 913
rect 44 807 78 841
rect 44 735 78 769
rect 44 663 78 697
rect 44 591 78 625
rect 44 519 78 553
rect 44 447 78 481
rect 44 375 78 409
rect 44 303 78 337
rect 44 231 78 265
rect 44 159 78 193
rect 44 87 78 121
rect 130 951 164 985
rect 130 879 164 913
rect 130 807 164 841
rect 130 735 164 769
rect 130 663 164 697
rect 130 591 164 625
rect 130 519 164 553
rect 130 447 164 481
rect 130 375 164 409
rect 130 303 164 337
rect 130 231 164 265
rect 130 159 164 193
rect 130 87 164 121
rect 216 951 250 985
rect 216 879 250 913
rect 216 807 250 841
rect 216 735 250 769
rect 216 663 250 697
rect 216 591 250 625
rect 216 519 250 553
rect 216 447 250 481
rect 216 375 250 409
rect 216 303 250 337
rect 216 231 250 265
rect 216 159 250 193
rect 216 87 250 121
<< poly >>
rect 80 1118 214 1134
rect 80 1084 96 1118
rect 130 1084 164 1118
rect 198 1084 214 1118
rect 80 1068 214 1084
rect 89 1062 205 1068
rect 89 1036 119 1062
rect 175 1036 205 1062
rect 89 10 119 36
rect 175 10 205 36
<< polycont >>
rect 96 1084 130 1118
rect 164 1084 198 1118
<< locali >>
rect 80 1118 214 1134
rect 80 1084 94 1118
rect 130 1084 164 1118
rect 200 1084 214 1118
rect 80 1068 214 1084
rect 44 985 78 1034
rect 44 913 78 951
rect 44 841 78 879
rect 44 769 78 807
rect 44 697 78 735
rect 44 625 78 663
rect 44 553 78 591
rect 44 481 78 519
rect 44 409 78 447
rect 44 337 78 375
rect 44 265 78 303
rect 44 193 78 231
rect 44 121 78 159
rect 44 36 78 87
rect 130 985 164 1034
rect 130 913 164 951
rect 130 841 164 879
rect 130 769 164 807
rect 130 697 164 735
rect 130 625 164 663
rect 130 553 164 591
rect 130 481 164 519
rect 130 409 164 447
rect 130 337 164 375
rect 130 265 164 303
rect 130 193 164 231
rect 130 121 164 159
rect 130 36 164 87
rect 216 985 250 1034
rect 216 913 250 951
rect 216 841 250 879
rect 216 769 250 807
rect 216 697 250 735
rect 216 625 250 663
rect 216 553 250 591
rect 216 481 250 519
rect 216 409 250 447
rect 216 337 250 375
rect 216 265 250 303
rect 216 193 250 231
rect 216 121 250 159
rect 216 36 250 87
<< viali >>
rect 94 1084 96 1118
rect 96 1084 128 1118
rect 166 1084 198 1118
rect 198 1084 200 1118
rect 44 951 78 985
rect 44 879 78 913
rect 44 807 78 841
rect 44 735 78 769
rect 44 663 78 697
rect 44 591 78 625
rect 44 519 78 553
rect 44 447 78 481
rect 44 375 78 409
rect 44 303 78 337
rect 44 231 78 265
rect 44 159 78 193
rect 44 87 78 121
rect 130 951 164 985
rect 130 879 164 913
rect 130 807 164 841
rect 130 735 164 769
rect 130 663 164 697
rect 130 591 164 625
rect 130 519 164 553
rect 130 447 164 481
rect 130 375 164 409
rect 130 303 164 337
rect 130 231 164 265
rect 130 159 164 193
rect 130 87 164 121
rect 216 951 250 985
rect 216 879 250 913
rect 216 807 250 841
rect 216 735 250 769
rect 216 663 250 697
rect 216 591 250 625
rect 216 519 250 553
rect 216 447 250 481
rect 216 375 250 409
rect 216 303 250 337
rect 216 231 250 265
rect 216 159 250 193
rect 216 87 250 121
<< metal1 >>
rect 82 1118 212 1130
rect 82 1084 94 1118
rect 128 1084 166 1118
rect 200 1084 212 1118
rect 82 1072 212 1084
rect 38 985 84 1034
rect 38 951 44 985
rect 78 951 84 985
rect 38 913 84 951
rect 38 879 44 913
rect 78 879 84 913
rect 38 841 84 879
rect 38 807 44 841
rect 78 807 84 841
rect 38 769 84 807
rect 38 735 44 769
rect 78 735 84 769
rect 38 697 84 735
rect 38 663 44 697
rect 78 663 84 697
rect 38 625 84 663
rect 38 591 44 625
rect 78 591 84 625
rect 38 553 84 591
rect 38 519 44 553
rect 78 519 84 553
rect 38 481 84 519
rect 38 447 44 481
rect 78 447 84 481
rect 38 409 84 447
rect 38 375 44 409
rect 78 375 84 409
rect 38 337 84 375
rect 38 303 44 337
rect 78 303 84 337
rect 38 265 84 303
rect 38 231 44 265
rect 78 231 84 265
rect 38 193 84 231
rect 38 159 44 193
rect 78 159 84 193
rect 38 121 84 159
rect 38 87 44 121
rect 78 87 84 121
rect 38 -45 84 87
rect 121 1026 173 1034
rect 121 962 130 974
rect 164 962 173 974
rect 121 879 130 910
rect 164 879 173 910
rect 121 841 173 879
rect 121 807 130 841
rect 164 807 173 841
rect 121 769 173 807
rect 121 735 130 769
rect 164 735 173 769
rect 121 697 173 735
rect 121 663 130 697
rect 164 663 173 697
rect 121 625 173 663
rect 121 591 130 625
rect 164 591 173 625
rect 121 553 173 591
rect 121 519 130 553
rect 164 519 173 553
rect 121 481 173 519
rect 121 447 130 481
rect 164 447 173 481
rect 121 409 173 447
rect 121 375 130 409
rect 164 375 173 409
rect 121 337 173 375
rect 121 303 130 337
rect 164 303 173 337
rect 121 265 173 303
rect 121 231 130 265
rect 164 231 173 265
rect 121 193 173 231
rect 121 159 130 193
rect 164 159 173 193
rect 121 121 173 159
rect 121 87 130 121
rect 164 87 173 121
rect 121 36 173 87
rect 210 985 256 1034
rect 210 951 216 985
rect 250 951 256 985
rect 210 913 256 951
rect 210 879 216 913
rect 250 879 256 913
rect 210 841 256 879
rect 210 807 216 841
rect 250 807 256 841
rect 210 769 256 807
rect 210 735 216 769
rect 250 735 256 769
rect 210 697 256 735
rect 210 663 216 697
rect 250 663 256 697
rect 210 625 256 663
rect 210 591 216 625
rect 250 591 256 625
rect 210 553 256 591
rect 210 519 216 553
rect 250 519 256 553
rect 210 481 256 519
rect 210 447 216 481
rect 250 447 256 481
rect 210 409 256 447
rect 210 375 216 409
rect 250 375 256 409
rect 210 337 256 375
rect 210 303 216 337
rect 250 303 256 337
rect 210 265 256 303
rect 210 231 216 265
rect 250 231 256 265
rect 210 193 256 231
rect 210 159 216 193
rect 250 159 256 193
rect 210 121 256 159
rect 210 87 216 121
rect 250 87 256 121
rect 210 -45 256 87
rect 38 -97 256 -45
<< via1 >>
rect 121 985 173 1026
rect 121 974 130 985
rect 130 974 164 985
rect 164 974 173 985
rect 121 951 130 962
rect 130 951 164 962
rect 164 951 173 962
rect 121 913 173 951
rect 121 910 130 913
rect 130 910 164 913
rect 164 910 173 913
<< metal2 >>
rect 121 1026 173 1032
rect 121 962 173 974
rect 121 904 173 910
<< labels >>
flabel metal2 s 121 904 173 1032 0 FreeSans 400 0 0 0 DRAIN
port 2 nsew
flabel metal1 s 38 -97 256 -45 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel metal1 s 82 1072 212 1130 0 FreeSans 400 0 0 0 GATE
port 4 nsew
flabel nwell s 74 1063 78 1070 0 FreeSans 400 0 0 0 BULK
port 5 nsew
<< properties >>
string GDS_END 10497040
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10488604
string path 1.525 25.850 1.525 -2.425 
<< end >>
