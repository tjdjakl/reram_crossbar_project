magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< dnwell >>
tri -700 6714 -614 6800 se
rect -614 6714 914 6800
tri 914 6714 1000 6800 sw
rect -700 -714 1000 6714
tri -700 -800 -614 -714 ne
rect -614 -800 914 -714
tri 914 -800 1000 -714 nw
<< nwell >>
rect -480 -560 780 6560
<< pwell >>
rect -1234 7074 1534 7208
rect -1234 6026 -1100 7074
rect -1234 -26 -574 6026
rect -1234 -1074 -1100 -26
rect 1400 6026 1534 7074
rect 874 -26 1534 6026
rect 1400 -1074 1534 -26
rect -1234 -1208 1534 -1074
<< mvnmos >>
rect -900 0 -730 6000
rect 1030 0 1200 6000
<< mvnnmos >>
rect -730 0 -600 6000
rect 900 0 1030 6000
<< mvndiff >>
rect -1026 5975 -900 6000
rect -1026 25 -1014 5975
rect -912 25 -900 5975
rect -1026 0 -900 25
rect 1200 5975 1326 6000
rect 1200 25 1212 5975
rect 1314 25 1326 5975
rect 1200 0 1326 25
<< mvndiffc >>
rect -1014 25 -912 5975
rect 1212 25 1314 5975
<< mvpsubdiff >>
rect -1208 7158 1508 7182
rect -1208 7124 -1159 7158
rect -1125 7124 -1091 7158
rect -1057 7124 -1023 7158
rect -989 7124 -955 7158
rect -921 7124 -887 7158
rect -853 7124 -819 7158
rect -785 7124 -751 7158
rect -717 7124 -683 7158
rect -649 7124 -615 7158
rect -581 7124 -547 7158
rect -513 7124 -479 7158
rect -445 7124 -411 7158
rect -377 7124 -343 7158
rect -309 7124 -275 7158
rect -241 7124 -207 7158
rect -173 7124 -139 7158
rect -105 7124 -71 7158
rect -37 7124 -3 7158
rect 31 7124 65 7158
rect 99 7124 133 7158
rect 167 7124 201 7158
rect 235 7124 269 7158
rect 303 7124 337 7158
rect 371 7124 405 7158
rect 439 7124 473 7158
rect 507 7124 541 7158
rect 575 7124 609 7158
rect 643 7124 677 7158
rect 711 7124 745 7158
rect 779 7124 813 7158
rect 847 7124 881 7158
rect 915 7124 949 7158
rect 983 7124 1017 7158
rect 1051 7124 1085 7158
rect 1119 7124 1153 7158
rect 1187 7124 1221 7158
rect 1255 7124 1289 7158
rect 1323 7124 1357 7158
rect 1391 7124 1425 7158
rect 1459 7124 1508 7158
rect -1208 7100 1508 7124
rect -1208 7063 -1126 7100
rect -1208 7029 -1184 7063
rect -1150 7029 -1126 7063
rect -1208 6995 -1126 7029
rect 1426 7063 1508 7100
rect 1426 7029 1450 7063
rect 1484 7029 1508 7063
rect -1208 6961 -1184 6995
rect -1150 6961 -1126 6995
rect -1208 6927 -1126 6961
rect -1208 6893 -1184 6927
rect -1150 6893 -1126 6927
rect -1208 6859 -1126 6893
rect -1208 6825 -1184 6859
rect -1150 6825 -1126 6859
rect -1208 6791 -1126 6825
rect -1208 6757 -1184 6791
rect -1150 6757 -1126 6791
rect -1208 6723 -1126 6757
rect -1208 6689 -1184 6723
rect -1150 6689 -1126 6723
rect -1208 6655 -1126 6689
rect -1208 6621 -1184 6655
rect -1150 6621 -1126 6655
rect -1208 6587 -1126 6621
rect -1208 6553 -1184 6587
rect -1150 6553 -1126 6587
rect -1208 6519 -1126 6553
rect -1208 6485 -1184 6519
rect -1150 6485 -1126 6519
rect -1208 6451 -1126 6485
rect -1208 6417 -1184 6451
rect -1150 6417 -1126 6451
rect -1208 6383 -1126 6417
rect -1208 6349 -1184 6383
rect -1150 6349 -1126 6383
rect -1208 6315 -1126 6349
rect -1208 6281 -1184 6315
rect -1150 6281 -1126 6315
rect -1208 6247 -1126 6281
rect -1208 6213 -1184 6247
rect -1150 6213 -1126 6247
rect -1208 6179 -1126 6213
rect -1208 6145 -1184 6179
rect -1150 6145 -1126 6179
rect -1208 6111 -1126 6145
rect -1208 6077 -1184 6111
rect -1150 6077 -1126 6111
rect -1208 6043 -1126 6077
rect -1208 6009 -1184 6043
rect -1150 6009 -1126 6043
rect -1208 5975 -1126 6009
rect 1426 6995 1508 7029
rect 1426 6961 1450 6995
rect 1484 6961 1508 6995
rect 1426 6927 1508 6961
rect 1426 6893 1450 6927
rect 1484 6893 1508 6927
rect 1426 6859 1508 6893
rect 1426 6825 1450 6859
rect 1484 6825 1508 6859
rect 1426 6791 1508 6825
rect 1426 6757 1450 6791
rect 1484 6757 1508 6791
rect 1426 6723 1508 6757
rect 1426 6689 1450 6723
rect 1484 6689 1508 6723
rect 1426 6655 1508 6689
rect 1426 6621 1450 6655
rect 1484 6621 1508 6655
rect 1426 6587 1508 6621
rect 1426 6553 1450 6587
rect 1484 6553 1508 6587
rect 1426 6519 1508 6553
rect 1426 6485 1450 6519
rect 1484 6485 1508 6519
rect 1426 6451 1508 6485
rect 1426 6417 1450 6451
rect 1484 6417 1508 6451
rect 1426 6383 1508 6417
rect 1426 6349 1450 6383
rect 1484 6349 1508 6383
rect 1426 6315 1508 6349
rect 1426 6281 1450 6315
rect 1484 6281 1508 6315
rect 1426 6247 1508 6281
rect 1426 6213 1450 6247
rect 1484 6213 1508 6247
rect 1426 6179 1508 6213
rect 1426 6145 1450 6179
rect 1484 6145 1508 6179
rect 1426 6111 1508 6145
rect 1426 6077 1450 6111
rect 1484 6077 1508 6111
rect 1426 6043 1508 6077
rect 1426 6009 1450 6043
rect 1484 6009 1508 6043
rect -1208 5941 -1184 5975
rect -1150 5941 -1126 5975
rect -1208 5907 -1126 5941
rect -1208 5873 -1184 5907
rect -1150 5873 -1126 5907
rect -1208 5839 -1126 5873
rect -1208 5805 -1184 5839
rect -1150 5805 -1126 5839
rect -1208 5771 -1126 5805
rect -1208 5737 -1184 5771
rect -1150 5737 -1126 5771
rect -1208 5703 -1126 5737
rect -1208 5669 -1184 5703
rect -1150 5669 -1126 5703
rect -1208 5635 -1126 5669
rect -1208 5601 -1184 5635
rect -1150 5601 -1126 5635
rect -1208 5567 -1126 5601
rect -1208 5533 -1184 5567
rect -1150 5533 -1126 5567
rect -1208 5499 -1126 5533
rect -1208 5465 -1184 5499
rect -1150 5465 -1126 5499
rect -1208 5431 -1126 5465
rect -1208 5397 -1184 5431
rect -1150 5397 -1126 5431
rect -1208 5363 -1126 5397
rect -1208 5329 -1184 5363
rect -1150 5329 -1126 5363
rect -1208 5295 -1126 5329
rect -1208 5261 -1184 5295
rect -1150 5261 -1126 5295
rect -1208 5227 -1126 5261
rect -1208 5193 -1184 5227
rect -1150 5193 -1126 5227
rect -1208 5159 -1126 5193
rect -1208 5125 -1184 5159
rect -1150 5125 -1126 5159
rect -1208 5091 -1126 5125
rect -1208 5057 -1184 5091
rect -1150 5057 -1126 5091
rect -1208 5023 -1126 5057
rect -1208 4989 -1184 5023
rect -1150 4989 -1126 5023
rect -1208 4955 -1126 4989
rect -1208 4921 -1184 4955
rect -1150 4921 -1126 4955
rect -1208 4887 -1126 4921
rect -1208 4853 -1184 4887
rect -1150 4853 -1126 4887
rect -1208 4819 -1126 4853
rect -1208 4785 -1184 4819
rect -1150 4785 -1126 4819
rect -1208 4751 -1126 4785
rect -1208 4717 -1184 4751
rect -1150 4717 -1126 4751
rect -1208 4683 -1126 4717
rect -1208 4649 -1184 4683
rect -1150 4649 -1126 4683
rect -1208 4615 -1126 4649
rect -1208 4581 -1184 4615
rect -1150 4581 -1126 4615
rect -1208 4547 -1126 4581
rect -1208 4513 -1184 4547
rect -1150 4513 -1126 4547
rect -1208 4479 -1126 4513
rect -1208 4445 -1184 4479
rect -1150 4445 -1126 4479
rect -1208 4411 -1126 4445
rect -1208 4377 -1184 4411
rect -1150 4377 -1126 4411
rect -1208 4343 -1126 4377
rect -1208 4309 -1184 4343
rect -1150 4309 -1126 4343
rect -1208 4275 -1126 4309
rect -1208 4241 -1184 4275
rect -1150 4241 -1126 4275
rect -1208 4207 -1126 4241
rect -1208 4173 -1184 4207
rect -1150 4173 -1126 4207
rect -1208 4139 -1126 4173
rect -1208 4105 -1184 4139
rect -1150 4105 -1126 4139
rect -1208 4071 -1126 4105
rect -1208 4037 -1184 4071
rect -1150 4037 -1126 4071
rect -1208 4003 -1126 4037
rect -1208 3969 -1184 4003
rect -1150 3969 -1126 4003
rect -1208 3935 -1126 3969
rect -1208 3901 -1184 3935
rect -1150 3901 -1126 3935
rect -1208 3867 -1126 3901
rect -1208 3833 -1184 3867
rect -1150 3833 -1126 3867
rect -1208 3799 -1126 3833
rect -1208 3765 -1184 3799
rect -1150 3765 -1126 3799
rect -1208 3731 -1126 3765
rect -1208 3697 -1184 3731
rect -1150 3697 -1126 3731
rect -1208 3663 -1126 3697
rect -1208 3629 -1184 3663
rect -1150 3629 -1126 3663
rect -1208 3595 -1126 3629
rect -1208 3561 -1184 3595
rect -1150 3561 -1126 3595
rect -1208 3527 -1126 3561
rect -1208 3493 -1184 3527
rect -1150 3493 -1126 3527
rect -1208 3459 -1126 3493
rect -1208 3425 -1184 3459
rect -1150 3425 -1126 3459
rect -1208 3391 -1126 3425
rect -1208 3357 -1184 3391
rect -1150 3357 -1126 3391
rect -1208 3323 -1126 3357
rect -1208 3289 -1184 3323
rect -1150 3289 -1126 3323
rect -1208 3255 -1126 3289
rect -1208 3221 -1184 3255
rect -1150 3221 -1126 3255
rect -1208 3187 -1126 3221
rect -1208 3153 -1184 3187
rect -1150 3153 -1126 3187
rect -1208 3119 -1126 3153
rect -1208 3085 -1184 3119
rect -1150 3085 -1126 3119
rect -1208 3051 -1126 3085
rect -1208 3017 -1184 3051
rect -1150 3017 -1126 3051
rect -1208 2983 -1126 3017
rect -1208 2949 -1184 2983
rect -1150 2949 -1126 2983
rect -1208 2915 -1126 2949
rect -1208 2881 -1184 2915
rect -1150 2881 -1126 2915
rect -1208 2847 -1126 2881
rect -1208 2813 -1184 2847
rect -1150 2813 -1126 2847
rect -1208 2779 -1126 2813
rect -1208 2745 -1184 2779
rect -1150 2745 -1126 2779
rect -1208 2711 -1126 2745
rect -1208 2677 -1184 2711
rect -1150 2677 -1126 2711
rect -1208 2643 -1126 2677
rect -1208 2609 -1184 2643
rect -1150 2609 -1126 2643
rect -1208 2575 -1126 2609
rect -1208 2541 -1184 2575
rect -1150 2541 -1126 2575
rect -1208 2507 -1126 2541
rect -1208 2473 -1184 2507
rect -1150 2473 -1126 2507
rect -1208 2439 -1126 2473
rect -1208 2405 -1184 2439
rect -1150 2405 -1126 2439
rect -1208 2371 -1126 2405
rect -1208 2337 -1184 2371
rect -1150 2337 -1126 2371
rect -1208 2303 -1126 2337
rect -1208 2269 -1184 2303
rect -1150 2269 -1126 2303
rect -1208 2235 -1126 2269
rect -1208 2201 -1184 2235
rect -1150 2201 -1126 2235
rect -1208 2167 -1126 2201
rect -1208 2133 -1184 2167
rect -1150 2133 -1126 2167
rect -1208 2099 -1126 2133
rect -1208 2065 -1184 2099
rect -1150 2065 -1126 2099
rect -1208 2031 -1126 2065
rect -1208 1997 -1184 2031
rect -1150 1997 -1126 2031
rect -1208 1963 -1126 1997
rect -1208 1929 -1184 1963
rect -1150 1929 -1126 1963
rect -1208 1895 -1126 1929
rect -1208 1861 -1184 1895
rect -1150 1861 -1126 1895
rect -1208 1827 -1126 1861
rect -1208 1793 -1184 1827
rect -1150 1793 -1126 1827
rect -1208 1759 -1126 1793
rect -1208 1725 -1184 1759
rect -1150 1725 -1126 1759
rect -1208 1691 -1126 1725
rect -1208 1657 -1184 1691
rect -1150 1657 -1126 1691
rect -1208 1623 -1126 1657
rect -1208 1589 -1184 1623
rect -1150 1589 -1126 1623
rect -1208 1555 -1126 1589
rect -1208 1521 -1184 1555
rect -1150 1521 -1126 1555
rect -1208 1487 -1126 1521
rect -1208 1453 -1184 1487
rect -1150 1453 -1126 1487
rect -1208 1419 -1126 1453
rect -1208 1385 -1184 1419
rect -1150 1385 -1126 1419
rect -1208 1351 -1126 1385
rect -1208 1317 -1184 1351
rect -1150 1317 -1126 1351
rect -1208 1283 -1126 1317
rect -1208 1249 -1184 1283
rect -1150 1249 -1126 1283
rect -1208 1215 -1126 1249
rect -1208 1181 -1184 1215
rect -1150 1181 -1126 1215
rect -1208 1147 -1126 1181
rect -1208 1113 -1184 1147
rect -1150 1113 -1126 1147
rect -1208 1079 -1126 1113
rect -1208 1045 -1184 1079
rect -1150 1045 -1126 1079
rect -1208 1011 -1126 1045
rect -1208 977 -1184 1011
rect -1150 977 -1126 1011
rect -1208 943 -1126 977
rect -1208 909 -1184 943
rect -1150 909 -1126 943
rect -1208 875 -1126 909
rect -1208 841 -1184 875
rect -1150 841 -1126 875
rect -1208 807 -1126 841
rect -1208 773 -1184 807
rect -1150 773 -1126 807
rect -1208 739 -1126 773
rect -1208 705 -1184 739
rect -1150 705 -1126 739
rect -1208 671 -1126 705
rect -1208 637 -1184 671
rect -1150 637 -1126 671
rect -1208 603 -1126 637
rect -1208 569 -1184 603
rect -1150 569 -1126 603
rect -1208 535 -1126 569
rect -1208 501 -1184 535
rect -1150 501 -1126 535
rect -1208 467 -1126 501
rect -1208 433 -1184 467
rect -1150 433 -1126 467
rect -1208 399 -1126 433
rect -1208 365 -1184 399
rect -1150 365 -1126 399
rect -1208 331 -1126 365
rect -1208 297 -1184 331
rect -1150 297 -1126 331
rect -1208 263 -1126 297
rect -1208 229 -1184 263
rect -1150 229 -1126 263
rect -1208 195 -1126 229
rect -1208 161 -1184 195
rect -1150 161 -1126 195
rect -1208 127 -1126 161
rect -1208 93 -1184 127
rect -1150 93 -1126 127
rect -1208 59 -1126 93
rect -1208 25 -1184 59
rect -1150 25 -1126 59
rect -1208 -9 -1126 25
rect 1426 5975 1508 6009
rect 1426 5941 1450 5975
rect 1484 5941 1508 5975
rect 1426 5907 1508 5941
rect 1426 5873 1450 5907
rect 1484 5873 1508 5907
rect 1426 5839 1508 5873
rect 1426 5805 1450 5839
rect 1484 5805 1508 5839
rect 1426 5771 1508 5805
rect 1426 5737 1450 5771
rect 1484 5737 1508 5771
rect 1426 5703 1508 5737
rect 1426 5669 1450 5703
rect 1484 5669 1508 5703
rect 1426 5635 1508 5669
rect 1426 5601 1450 5635
rect 1484 5601 1508 5635
rect 1426 5567 1508 5601
rect 1426 5533 1450 5567
rect 1484 5533 1508 5567
rect 1426 5499 1508 5533
rect 1426 5465 1450 5499
rect 1484 5465 1508 5499
rect 1426 5431 1508 5465
rect 1426 5397 1450 5431
rect 1484 5397 1508 5431
rect 1426 5363 1508 5397
rect 1426 5329 1450 5363
rect 1484 5329 1508 5363
rect 1426 5295 1508 5329
rect 1426 5261 1450 5295
rect 1484 5261 1508 5295
rect 1426 5227 1508 5261
rect 1426 5193 1450 5227
rect 1484 5193 1508 5227
rect 1426 5159 1508 5193
rect 1426 5125 1450 5159
rect 1484 5125 1508 5159
rect 1426 5091 1508 5125
rect 1426 5057 1450 5091
rect 1484 5057 1508 5091
rect 1426 5023 1508 5057
rect 1426 4989 1450 5023
rect 1484 4989 1508 5023
rect 1426 4955 1508 4989
rect 1426 4921 1450 4955
rect 1484 4921 1508 4955
rect 1426 4887 1508 4921
rect 1426 4853 1450 4887
rect 1484 4853 1508 4887
rect 1426 4819 1508 4853
rect 1426 4785 1450 4819
rect 1484 4785 1508 4819
rect 1426 4751 1508 4785
rect 1426 4717 1450 4751
rect 1484 4717 1508 4751
rect 1426 4683 1508 4717
rect 1426 4649 1450 4683
rect 1484 4649 1508 4683
rect 1426 4615 1508 4649
rect 1426 4581 1450 4615
rect 1484 4581 1508 4615
rect 1426 4547 1508 4581
rect 1426 4513 1450 4547
rect 1484 4513 1508 4547
rect 1426 4479 1508 4513
rect 1426 4445 1450 4479
rect 1484 4445 1508 4479
rect 1426 4411 1508 4445
rect 1426 4377 1450 4411
rect 1484 4377 1508 4411
rect 1426 4343 1508 4377
rect 1426 4309 1450 4343
rect 1484 4309 1508 4343
rect 1426 4275 1508 4309
rect 1426 4241 1450 4275
rect 1484 4241 1508 4275
rect 1426 4207 1508 4241
rect 1426 4173 1450 4207
rect 1484 4173 1508 4207
rect 1426 4139 1508 4173
rect 1426 4105 1450 4139
rect 1484 4105 1508 4139
rect 1426 4071 1508 4105
rect 1426 4037 1450 4071
rect 1484 4037 1508 4071
rect 1426 4003 1508 4037
rect 1426 3969 1450 4003
rect 1484 3969 1508 4003
rect 1426 3935 1508 3969
rect 1426 3901 1450 3935
rect 1484 3901 1508 3935
rect 1426 3867 1508 3901
rect 1426 3833 1450 3867
rect 1484 3833 1508 3867
rect 1426 3799 1508 3833
rect 1426 3765 1450 3799
rect 1484 3765 1508 3799
rect 1426 3731 1508 3765
rect 1426 3697 1450 3731
rect 1484 3697 1508 3731
rect 1426 3663 1508 3697
rect 1426 3629 1450 3663
rect 1484 3629 1508 3663
rect 1426 3595 1508 3629
rect 1426 3561 1450 3595
rect 1484 3561 1508 3595
rect 1426 3527 1508 3561
rect 1426 3493 1450 3527
rect 1484 3493 1508 3527
rect 1426 3459 1508 3493
rect 1426 3425 1450 3459
rect 1484 3425 1508 3459
rect 1426 3391 1508 3425
rect 1426 3357 1450 3391
rect 1484 3357 1508 3391
rect 1426 3323 1508 3357
rect 1426 3289 1450 3323
rect 1484 3289 1508 3323
rect 1426 3255 1508 3289
rect 1426 3221 1450 3255
rect 1484 3221 1508 3255
rect 1426 3187 1508 3221
rect 1426 3153 1450 3187
rect 1484 3153 1508 3187
rect 1426 3119 1508 3153
rect 1426 3085 1450 3119
rect 1484 3085 1508 3119
rect 1426 3051 1508 3085
rect 1426 3017 1450 3051
rect 1484 3017 1508 3051
rect 1426 2983 1508 3017
rect 1426 2949 1450 2983
rect 1484 2949 1508 2983
rect 1426 2915 1508 2949
rect 1426 2881 1450 2915
rect 1484 2881 1508 2915
rect 1426 2847 1508 2881
rect 1426 2813 1450 2847
rect 1484 2813 1508 2847
rect 1426 2779 1508 2813
rect 1426 2745 1450 2779
rect 1484 2745 1508 2779
rect 1426 2711 1508 2745
rect 1426 2677 1450 2711
rect 1484 2677 1508 2711
rect 1426 2643 1508 2677
rect 1426 2609 1450 2643
rect 1484 2609 1508 2643
rect 1426 2575 1508 2609
rect 1426 2541 1450 2575
rect 1484 2541 1508 2575
rect 1426 2507 1508 2541
rect 1426 2473 1450 2507
rect 1484 2473 1508 2507
rect 1426 2439 1508 2473
rect 1426 2405 1450 2439
rect 1484 2405 1508 2439
rect 1426 2371 1508 2405
rect 1426 2337 1450 2371
rect 1484 2337 1508 2371
rect 1426 2303 1508 2337
rect 1426 2269 1450 2303
rect 1484 2269 1508 2303
rect 1426 2235 1508 2269
rect 1426 2201 1450 2235
rect 1484 2201 1508 2235
rect 1426 2167 1508 2201
rect 1426 2133 1450 2167
rect 1484 2133 1508 2167
rect 1426 2099 1508 2133
rect 1426 2065 1450 2099
rect 1484 2065 1508 2099
rect 1426 2031 1508 2065
rect 1426 1997 1450 2031
rect 1484 1997 1508 2031
rect 1426 1963 1508 1997
rect 1426 1929 1450 1963
rect 1484 1929 1508 1963
rect 1426 1895 1508 1929
rect 1426 1861 1450 1895
rect 1484 1861 1508 1895
rect 1426 1827 1508 1861
rect 1426 1793 1450 1827
rect 1484 1793 1508 1827
rect 1426 1759 1508 1793
rect 1426 1725 1450 1759
rect 1484 1725 1508 1759
rect 1426 1691 1508 1725
rect 1426 1657 1450 1691
rect 1484 1657 1508 1691
rect 1426 1623 1508 1657
rect 1426 1589 1450 1623
rect 1484 1589 1508 1623
rect 1426 1555 1508 1589
rect 1426 1521 1450 1555
rect 1484 1521 1508 1555
rect 1426 1487 1508 1521
rect 1426 1453 1450 1487
rect 1484 1453 1508 1487
rect 1426 1419 1508 1453
rect 1426 1385 1450 1419
rect 1484 1385 1508 1419
rect 1426 1351 1508 1385
rect 1426 1317 1450 1351
rect 1484 1317 1508 1351
rect 1426 1283 1508 1317
rect 1426 1249 1450 1283
rect 1484 1249 1508 1283
rect 1426 1215 1508 1249
rect 1426 1181 1450 1215
rect 1484 1181 1508 1215
rect 1426 1147 1508 1181
rect 1426 1113 1450 1147
rect 1484 1113 1508 1147
rect 1426 1079 1508 1113
rect 1426 1045 1450 1079
rect 1484 1045 1508 1079
rect 1426 1011 1508 1045
rect 1426 977 1450 1011
rect 1484 977 1508 1011
rect 1426 943 1508 977
rect 1426 909 1450 943
rect 1484 909 1508 943
rect 1426 875 1508 909
rect 1426 841 1450 875
rect 1484 841 1508 875
rect 1426 807 1508 841
rect 1426 773 1450 807
rect 1484 773 1508 807
rect 1426 739 1508 773
rect 1426 705 1450 739
rect 1484 705 1508 739
rect 1426 671 1508 705
rect 1426 637 1450 671
rect 1484 637 1508 671
rect 1426 603 1508 637
rect 1426 569 1450 603
rect 1484 569 1508 603
rect 1426 535 1508 569
rect 1426 501 1450 535
rect 1484 501 1508 535
rect 1426 467 1508 501
rect 1426 433 1450 467
rect 1484 433 1508 467
rect 1426 399 1508 433
rect 1426 365 1450 399
rect 1484 365 1508 399
rect 1426 331 1508 365
rect 1426 297 1450 331
rect 1484 297 1508 331
rect 1426 263 1508 297
rect 1426 229 1450 263
rect 1484 229 1508 263
rect 1426 195 1508 229
rect 1426 161 1450 195
rect 1484 161 1508 195
rect 1426 127 1508 161
rect 1426 93 1450 127
rect 1484 93 1508 127
rect 1426 59 1508 93
rect 1426 25 1450 59
rect 1484 25 1508 59
rect -1208 -43 -1184 -9
rect -1150 -43 -1126 -9
rect -1208 -77 -1126 -43
rect -1208 -111 -1184 -77
rect -1150 -111 -1126 -77
rect -1208 -145 -1126 -111
rect -1208 -179 -1184 -145
rect -1150 -179 -1126 -145
rect -1208 -213 -1126 -179
rect -1208 -247 -1184 -213
rect -1150 -247 -1126 -213
rect -1208 -281 -1126 -247
rect -1208 -315 -1184 -281
rect -1150 -315 -1126 -281
rect -1208 -349 -1126 -315
rect -1208 -383 -1184 -349
rect -1150 -383 -1126 -349
rect -1208 -417 -1126 -383
rect -1208 -451 -1184 -417
rect -1150 -451 -1126 -417
rect -1208 -485 -1126 -451
rect -1208 -519 -1184 -485
rect -1150 -519 -1126 -485
rect -1208 -553 -1126 -519
rect -1208 -587 -1184 -553
rect -1150 -587 -1126 -553
rect -1208 -621 -1126 -587
rect -1208 -655 -1184 -621
rect -1150 -655 -1126 -621
rect -1208 -689 -1126 -655
rect -1208 -723 -1184 -689
rect -1150 -723 -1126 -689
rect -1208 -757 -1126 -723
rect -1208 -791 -1184 -757
rect -1150 -791 -1126 -757
rect -1208 -825 -1126 -791
rect -1208 -859 -1184 -825
rect -1150 -859 -1126 -825
rect -1208 -893 -1126 -859
rect -1208 -927 -1184 -893
rect -1150 -927 -1126 -893
rect -1208 -961 -1126 -927
rect -1208 -995 -1184 -961
rect -1150 -995 -1126 -961
rect -1208 -1029 -1126 -995
rect 1426 -9 1508 25
rect 1426 -43 1450 -9
rect 1484 -43 1508 -9
rect 1426 -77 1508 -43
rect 1426 -111 1450 -77
rect 1484 -111 1508 -77
rect 1426 -145 1508 -111
rect 1426 -179 1450 -145
rect 1484 -179 1508 -145
rect 1426 -213 1508 -179
rect 1426 -247 1450 -213
rect 1484 -247 1508 -213
rect 1426 -281 1508 -247
rect 1426 -315 1450 -281
rect 1484 -315 1508 -281
rect 1426 -349 1508 -315
rect 1426 -383 1450 -349
rect 1484 -383 1508 -349
rect 1426 -417 1508 -383
rect 1426 -451 1450 -417
rect 1484 -451 1508 -417
rect 1426 -485 1508 -451
rect 1426 -519 1450 -485
rect 1484 -519 1508 -485
rect 1426 -553 1508 -519
rect 1426 -587 1450 -553
rect 1484 -587 1508 -553
rect 1426 -621 1508 -587
rect 1426 -655 1450 -621
rect 1484 -655 1508 -621
rect 1426 -689 1508 -655
rect 1426 -723 1450 -689
rect 1484 -723 1508 -689
rect 1426 -757 1508 -723
rect 1426 -791 1450 -757
rect 1484 -791 1508 -757
rect 1426 -825 1508 -791
rect 1426 -859 1450 -825
rect 1484 -859 1508 -825
rect 1426 -893 1508 -859
rect 1426 -927 1450 -893
rect 1484 -927 1508 -893
rect 1426 -961 1508 -927
rect 1426 -995 1450 -961
rect 1484 -995 1508 -961
rect -1208 -1063 -1184 -1029
rect -1150 -1063 -1126 -1029
rect -1208 -1100 -1126 -1063
rect 1426 -1029 1508 -995
rect 1426 -1063 1450 -1029
rect 1484 -1063 1508 -1029
rect 1426 -1100 1508 -1063
rect -1208 -1124 1508 -1100
rect -1208 -1158 -1159 -1124
rect -1125 -1158 -1091 -1124
rect -1057 -1158 -1023 -1124
rect -989 -1158 -955 -1124
rect -921 -1158 -887 -1124
rect -853 -1158 -819 -1124
rect -785 -1158 -751 -1124
rect -717 -1158 -683 -1124
rect -649 -1158 -615 -1124
rect -581 -1158 -547 -1124
rect -513 -1158 -479 -1124
rect -445 -1158 -411 -1124
rect -377 -1158 -343 -1124
rect -309 -1158 -275 -1124
rect -241 -1158 -207 -1124
rect -173 -1158 -139 -1124
rect -105 -1158 -71 -1124
rect -37 -1158 -3 -1124
rect 31 -1158 65 -1124
rect 99 -1158 133 -1124
rect 167 -1158 201 -1124
rect 235 -1158 269 -1124
rect 303 -1158 337 -1124
rect 371 -1158 405 -1124
rect 439 -1158 473 -1124
rect 507 -1158 541 -1124
rect 575 -1158 609 -1124
rect 643 -1158 677 -1124
rect 711 -1158 745 -1124
rect 779 -1158 813 -1124
rect 847 -1158 881 -1124
rect 915 -1158 949 -1124
rect 983 -1158 1017 -1124
rect 1051 -1158 1085 -1124
rect 1119 -1158 1153 -1124
rect 1187 -1158 1221 -1124
rect 1255 -1158 1289 -1124
rect 1323 -1158 1357 -1124
rect 1391 -1158 1425 -1124
rect 1459 -1158 1508 -1124
rect -1208 -1182 1508 -1158
<< mvnsubdiff >>
tri 0 5970 30 6000 se
rect 30 5970 270 6000
tri 270 5970 300 6000 sw
rect 0 5941 300 5970
rect 0 59 31 5941
rect 269 59 300 5941
rect 0 30 300 59
tri 0 0 30 30 ne
rect 30 0 270 30
tri 270 0 300 30 nw
<< mvpsubdiffcont >>
rect -1159 7124 -1125 7158
rect -1091 7124 -1057 7158
rect -1023 7124 -989 7158
rect -955 7124 -921 7158
rect -887 7124 -853 7158
rect -819 7124 -785 7158
rect -751 7124 -717 7158
rect -683 7124 -649 7158
rect -615 7124 -581 7158
rect -547 7124 -513 7158
rect -479 7124 -445 7158
rect -411 7124 -377 7158
rect -343 7124 -309 7158
rect -275 7124 -241 7158
rect -207 7124 -173 7158
rect -139 7124 -105 7158
rect -71 7124 -37 7158
rect -3 7124 31 7158
rect 65 7124 99 7158
rect 133 7124 167 7158
rect 201 7124 235 7158
rect 269 7124 303 7158
rect 337 7124 371 7158
rect 405 7124 439 7158
rect 473 7124 507 7158
rect 541 7124 575 7158
rect 609 7124 643 7158
rect 677 7124 711 7158
rect 745 7124 779 7158
rect 813 7124 847 7158
rect 881 7124 915 7158
rect 949 7124 983 7158
rect 1017 7124 1051 7158
rect 1085 7124 1119 7158
rect 1153 7124 1187 7158
rect 1221 7124 1255 7158
rect 1289 7124 1323 7158
rect 1357 7124 1391 7158
rect 1425 7124 1459 7158
rect -1184 7029 -1150 7063
rect 1450 7029 1484 7063
rect -1184 6961 -1150 6995
rect -1184 6893 -1150 6927
rect -1184 6825 -1150 6859
rect -1184 6757 -1150 6791
rect -1184 6689 -1150 6723
rect -1184 6621 -1150 6655
rect -1184 6553 -1150 6587
rect -1184 6485 -1150 6519
rect -1184 6417 -1150 6451
rect -1184 6349 -1150 6383
rect -1184 6281 -1150 6315
rect -1184 6213 -1150 6247
rect -1184 6145 -1150 6179
rect -1184 6077 -1150 6111
rect -1184 6009 -1150 6043
rect 1450 6961 1484 6995
rect 1450 6893 1484 6927
rect 1450 6825 1484 6859
rect 1450 6757 1484 6791
rect 1450 6689 1484 6723
rect 1450 6621 1484 6655
rect 1450 6553 1484 6587
rect 1450 6485 1484 6519
rect 1450 6417 1484 6451
rect 1450 6349 1484 6383
rect 1450 6281 1484 6315
rect 1450 6213 1484 6247
rect 1450 6145 1484 6179
rect 1450 6077 1484 6111
rect 1450 6009 1484 6043
rect -1184 5941 -1150 5975
rect -1184 5873 -1150 5907
rect -1184 5805 -1150 5839
rect -1184 5737 -1150 5771
rect -1184 5669 -1150 5703
rect -1184 5601 -1150 5635
rect -1184 5533 -1150 5567
rect -1184 5465 -1150 5499
rect -1184 5397 -1150 5431
rect -1184 5329 -1150 5363
rect -1184 5261 -1150 5295
rect -1184 5193 -1150 5227
rect -1184 5125 -1150 5159
rect -1184 5057 -1150 5091
rect -1184 4989 -1150 5023
rect -1184 4921 -1150 4955
rect -1184 4853 -1150 4887
rect -1184 4785 -1150 4819
rect -1184 4717 -1150 4751
rect -1184 4649 -1150 4683
rect -1184 4581 -1150 4615
rect -1184 4513 -1150 4547
rect -1184 4445 -1150 4479
rect -1184 4377 -1150 4411
rect -1184 4309 -1150 4343
rect -1184 4241 -1150 4275
rect -1184 4173 -1150 4207
rect -1184 4105 -1150 4139
rect -1184 4037 -1150 4071
rect -1184 3969 -1150 4003
rect -1184 3901 -1150 3935
rect -1184 3833 -1150 3867
rect -1184 3765 -1150 3799
rect -1184 3697 -1150 3731
rect -1184 3629 -1150 3663
rect -1184 3561 -1150 3595
rect -1184 3493 -1150 3527
rect -1184 3425 -1150 3459
rect -1184 3357 -1150 3391
rect -1184 3289 -1150 3323
rect -1184 3221 -1150 3255
rect -1184 3153 -1150 3187
rect -1184 3085 -1150 3119
rect -1184 3017 -1150 3051
rect -1184 2949 -1150 2983
rect -1184 2881 -1150 2915
rect -1184 2813 -1150 2847
rect -1184 2745 -1150 2779
rect -1184 2677 -1150 2711
rect -1184 2609 -1150 2643
rect -1184 2541 -1150 2575
rect -1184 2473 -1150 2507
rect -1184 2405 -1150 2439
rect -1184 2337 -1150 2371
rect -1184 2269 -1150 2303
rect -1184 2201 -1150 2235
rect -1184 2133 -1150 2167
rect -1184 2065 -1150 2099
rect -1184 1997 -1150 2031
rect -1184 1929 -1150 1963
rect -1184 1861 -1150 1895
rect -1184 1793 -1150 1827
rect -1184 1725 -1150 1759
rect -1184 1657 -1150 1691
rect -1184 1589 -1150 1623
rect -1184 1521 -1150 1555
rect -1184 1453 -1150 1487
rect -1184 1385 -1150 1419
rect -1184 1317 -1150 1351
rect -1184 1249 -1150 1283
rect -1184 1181 -1150 1215
rect -1184 1113 -1150 1147
rect -1184 1045 -1150 1079
rect -1184 977 -1150 1011
rect -1184 909 -1150 943
rect -1184 841 -1150 875
rect -1184 773 -1150 807
rect -1184 705 -1150 739
rect -1184 637 -1150 671
rect -1184 569 -1150 603
rect -1184 501 -1150 535
rect -1184 433 -1150 467
rect -1184 365 -1150 399
rect -1184 297 -1150 331
rect -1184 229 -1150 263
rect -1184 161 -1150 195
rect -1184 93 -1150 127
rect -1184 25 -1150 59
rect 1450 5941 1484 5975
rect 1450 5873 1484 5907
rect 1450 5805 1484 5839
rect 1450 5737 1484 5771
rect 1450 5669 1484 5703
rect 1450 5601 1484 5635
rect 1450 5533 1484 5567
rect 1450 5465 1484 5499
rect 1450 5397 1484 5431
rect 1450 5329 1484 5363
rect 1450 5261 1484 5295
rect 1450 5193 1484 5227
rect 1450 5125 1484 5159
rect 1450 5057 1484 5091
rect 1450 4989 1484 5023
rect 1450 4921 1484 4955
rect 1450 4853 1484 4887
rect 1450 4785 1484 4819
rect 1450 4717 1484 4751
rect 1450 4649 1484 4683
rect 1450 4581 1484 4615
rect 1450 4513 1484 4547
rect 1450 4445 1484 4479
rect 1450 4377 1484 4411
rect 1450 4309 1484 4343
rect 1450 4241 1484 4275
rect 1450 4173 1484 4207
rect 1450 4105 1484 4139
rect 1450 4037 1484 4071
rect 1450 3969 1484 4003
rect 1450 3901 1484 3935
rect 1450 3833 1484 3867
rect 1450 3765 1484 3799
rect 1450 3697 1484 3731
rect 1450 3629 1484 3663
rect 1450 3561 1484 3595
rect 1450 3493 1484 3527
rect 1450 3425 1484 3459
rect 1450 3357 1484 3391
rect 1450 3289 1484 3323
rect 1450 3221 1484 3255
rect 1450 3153 1484 3187
rect 1450 3085 1484 3119
rect 1450 3017 1484 3051
rect 1450 2949 1484 2983
rect 1450 2881 1484 2915
rect 1450 2813 1484 2847
rect 1450 2745 1484 2779
rect 1450 2677 1484 2711
rect 1450 2609 1484 2643
rect 1450 2541 1484 2575
rect 1450 2473 1484 2507
rect 1450 2405 1484 2439
rect 1450 2337 1484 2371
rect 1450 2269 1484 2303
rect 1450 2201 1484 2235
rect 1450 2133 1484 2167
rect 1450 2065 1484 2099
rect 1450 1997 1484 2031
rect 1450 1929 1484 1963
rect 1450 1861 1484 1895
rect 1450 1793 1484 1827
rect 1450 1725 1484 1759
rect 1450 1657 1484 1691
rect 1450 1589 1484 1623
rect 1450 1521 1484 1555
rect 1450 1453 1484 1487
rect 1450 1385 1484 1419
rect 1450 1317 1484 1351
rect 1450 1249 1484 1283
rect 1450 1181 1484 1215
rect 1450 1113 1484 1147
rect 1450 1045 1484 1079
rect 1450 977 1484 1011
rect 1450 909 1484 943
rect 1450 841 1484 875
rect 1450 773 1484 807
rect 1450 705 1484 739
rect 1450 637 1484 671
rect 1450 569 1484 603
rect 1450 501 1484 535
rect 1450 433 1484 467
rect 1450 365 1484 399
rect 1450 297 1484 331
rect 1450 229 1484 263
rect 1450 161 1484 195
rect 1450 93 1484 127
rect 1450 25 1484 59
rect -1184 -43 -1150 -9
rect -1184 -111 -1150 -77
rect -1184 -179 -1150 -145
rect -1184 -247 -1150 -213
rect -1184 -315 -1150 -281
rect -1184 -383 -1150 -349
rect -1184 -451 -1150 -417
rect -1184 -519 -1150 -485
rect -1184 -587 -1150 -553
rect -1184 -655 -1150 -621
rect -1184 -723 -1150 -689
rect -1184 -791 -1150 -757
rect -1184 -859 -1150 -825
rect -1184 -927 -1150 -893
rect -1184 -995 -1150 -961
rect 1450 -43 1484 -9
rect 1450 -111 1484 -77
rect 1450 -179 1484 -145
rect 1450 -247 1484 -213
rect 1450 -315 1484 -281
rect 1450 -383 1484 -349
rect 1450 -451 1484 -417
rect 1450 -519 1484 -485
rect 1450 -587 1484 -553
rect 1450 -655 1484 -621
rect 1450 -723 1484 -689
rect 1450 -791 1484 -757
rect 1450 -859 1484 -825
rect 1450 -927 1484 -893
rect 1450 -995 1484 -961
rect -1184 -1063 -1150 -1029
rect 1450 -1063 1484 -1029
rect -1159 -1158 -1125 -1124
rect -1091 -1158 -1057 -1124
rect -1023 -1158 -989 -1124
rect -955 -1158 -921 -1124
rect -887 -1158 -853 -1124
rect -819 -1158 -785 -1124
rect -751 -1158 -717 -1124
rect -683 -1158 -649 -1124
rect -615 -1158 -581 -1124
rect -547 -1158 -513 -1124
rect -479 -1158 -445 -1124
rect -411 -1158 -377 -1124
rect -343 -1158 -309 -1124
rect -275 -1158 -241 -1124
rect -207 -1158 -173 -1124
rect -139 -1158 -105 -1124
rect -71 -1158 -37 -1124
rect -3 -1158 31 -1124
rect 65 -1158 99 -1124
rect 133 -1158 167 -1124
rect 201 -1158 235 -1124
rect 269 -1158 303 -1124
rect 337 -1158 371 -1124
rect 405 -1158 439 -1124
rect 473 -1158 507 -1124
rect 541 -1158 575 -1124
rect 609 -1158 643 -1124
rect 677 -1158 711 -1124
rect 745 -1158 779 -1124
rect 813 -1158 847 -1124
rect 881 -1158 915 -1124
rect 949 -1158 983 -1124
rect 1017 -1158 1051 -1124
rect 1085 -1158 1119 -1124
rect 1153 -1158 1187 -1124
rect 1221 -1158 1255 -1124
rect 1289 -1158 1323 -1124
rect 1357 -1158 1391 -1124
rect 1425 -1158 1459 -1124
<< mvnsubdiffcont >>
rect 31 59 269 5941
<< poly >>
rect -900 6400 1200 7000
rect -900 6000 -300 6400
rect 600 6000 1200 6400
rect -600 0 -300 6000
rect 600 0 900 6000
rect -900 -400 -300 0
rect 600 -400 1200 0
rect -900 -665 1200 -400
rect -900 -835 -173 -665
rect 473 -835 1200 -665
rect -900 -1000 1200 -835
<< polycont >>
rect -173 -835 473 -665
<< locali >>
rect -1208 7158 1508 7182
rect -1208 7157 -1159 7158
rect -1125 7157 -1091 7158
rect -1057 7157 -1023 7158
rect -989 7157 -955 7158
rect -921 7157 -887 7158
rect -1208 7063 -1162 7157
rect -912 7124 -887 7157
rect -853 7157 -819 7158
rect -785 7157 -751 7158
rect -717 7157 -683 7158
rect -649 7157 -615 7158
rect -581 7157 -547 7158
rect -513 7157 -479 7158
rect -445 7157 -411 7158
rect -377 7157 -343 7158
rect -309 7157 -275 7158
rect -241 7157 -207 7158
rect -173 7157 -139 7158
rect -105 7157 -71 7158
rect -37 7157 -3 7158
rect 31 7157 65 7158
rect 99 7157 133 7158
rect 167 7157 201 7158
rect 235 7157 269 7158
rect 303 7157 337 7158
rect 371 7157 405 7158
rect 439 7157 473 7158
rect 507 7157 541 7158
rect 575 7157 609 7158
rect 643 7157 677 7158
rect 711 7157 745 7158
rect 779 7157 813 7158
rect 847 7157 881 7158
rect 915 7157 949 7158
rect 983 7157 1017 7158
rect 1051 7157 1085 7158
rect 1119 7157 1153 7158
rect -853 7124 -839 7157
rect 1139 7124 1153 7157
rect 1187 7157 1221 7158
rect 1255 7157 1289 7158
rect 1323 7157 1357 7158
rect 1391 7157 1425 7158
rect 1459 7157 1508 7158
rect 1187 7124 1212 7157
rect -1208 7029 -1184 7063
rect -1208 6995 -1162 7029
rect -1208 6961 -1184 6995
rect -1208 6927 -1162 6961
rect -1208 6893 -1184 6927
rect -912 6907 -839 7124
rect 1139 6907 1212 7124
rect 1462 7063 1508 7157
rect 1484 7029 1508 7063
rect 1462 6995 1508 7029
rect 1484 6961 1508 6995
rect 1462 6927 1508 6961
rect -1208 6859 -1162 6893
rect -912 6870 1212 6907
rect 1484 6893 1508 6927
rect -1208 6825 -1184 6859
rect -1208 6791 -1162 6825
rect -1208 6757 -1184 6791
rect -1208 6723 -1162 6757
rect -1208 6689 -1184 6723
rect -1208 6655 -1162 6689
rect -1208 6621 -1184 6655
rect -1208 6587 -1162 6621
rect -1208 6553 -1184 6587
rect -1208 6519 -1162 6553
rect -1208 6485 -1184 6519
rect -1208 6451 -1162 6485
rect -1208 6417 -1184 6451
rect -1208 6383 -1162 6417
rect -1208 6349 -1184 6383
rect -1208 6315 -1162 6349
rect -1208 6281 -1184 6315
rect -1208 6247 -1162 6281
rect -1208 6213 -1184 6247
rect -1208 6179 -1162 6213
rect -1208 6145 -1184 6179
rect -1208 6111 -1162 6145
rect -1208 6077 -1184 6111
rect -1208 6043 -1162 6077
rect -1208 6009 -1184 6043
rect -1208 5975 -1162 6009
rect -1208 5941 -1184 5975
rect -1208 5907 -1162 5941
rect -1208 5873 -1184 5907
rect -1208 5839 -1162 5873
rect -1208 5805 -1184 5839
rect -1208 5771 -1162 5805
rect -1208 5737 -1184 5771
rect -1208 5703 -1162 5737
rect -1208 5669 -1184 5703
rect -1208 5635 -1162 5669
rect -1208 5601 -1184 5635
rect -1208 5567 -1162 5601
rect -1208 5533 -1184 5567
rect -1208 5499 -1162 5533
rect -1208 5465 -1184 5499
rect -1208 5431 -1162 5465
rect -1208 5397 -1184 5431
rect -1208 5363 -1162 5397
rect -1208 5329 -1184 5363
rect -1208 5295 -1162 5329
rect -1208 5261 -1184 5295
rect -1208 5227 -1162 5261
rect -1208 5193 -1184 5227
rect -1208 5159 -1162 5193
rect -1208 5125 -1184 5159
rect -1208 5091 -1162 5125
rect -1208 5057 -1184 5091
rect -1208 5023 -1162 5057
rect -1208 4989 -1184 5023
rect -1208 4955 -1162 4989
rect -1208 4921 -1184 4955
rect -1208 4887 -1162 4921
rect -1208 4853 -1184 4887
rect -1208 4819 -1162 4853
rect -1208 4785 -1184 4819
rect -1208 4751 -1162 4785
rect -1208 4717 -1184 4751
rect -1208 4683 -1162 4717
rect -1208 4649 -1184 4683
rect -1208 4615 -1162 4649
rect -1208 4581 -1184 4615
rect -1208 4547 -1162 4581
rect -1208 4513 -1184 4547
rect -1208 4479 -1162 4513
rect -1208 4445 -1184 4479
rect -1208 4411 -1162 4445
rect -1208 4377 -1184 4411
rect -1208 4343 -1162 4377
rect -1208 4309 -1184 4343
rect -1208 4275 -1162 4309
rect -1208 4241 -1184 4275
rect -1208 4207 -1162 4241
rect -1208 4173 -1184 4207
rect -1208 4139 -1162 4173
rect -1208 4105 -1184 4139
rect -1208 4071 -1162 4105
rect -1208 4037 -1184 4071
rect -1208 4003 -1162 4037
rect -1208 3969 -1184 4003
rect -1208 3935 -1162 3969
rect -1208 3901 -1184 3935
rect -1208 3867 -1162 3901
rect -1208 3833 -1184 3867
rect -1208 3799 -1162 3833
rect -1208 3765 -1184 3799
rect -1208 3731 -1162 3765
rect -1208 3697 -1184 3731
rect -1208 3663 -1162 3697
rect -1208 3629 -1184 3663
rect -1208 3595 -1162 3629
rect -1208 3561 -1184 3595
rect -1208 3527 -1162 3561
rect -1208 3493 -1184 3527
rect -1208 3459 -1162 3493
rect -1208 3425 -1184 3459
rect -1208 3391 -1162 3425
rect -1208 3357 -1184 3391
rect -1208 3323 -1162 3357
rect -1208 3289 -1184 3323
rect -1208 3255 -1162 3289
rect -1208 3221 -1184 3255
rect -1208 3187 -1162 3221
rect -1208 3153 -1184 3187
rect -1208 3119 -1162 3153
rect -1208 3085 -1184 3119
rect -1208 3051 -1162 3085
rect -1208 3017 -1184 3051
rect -1208 2983 -1162 3017
rect -1208 2949 -1184 2983
rect -1208 2915 -1162 2949
rect -1208 2881 -1184 2915
rect -1208 2847 -1162 2881
rect -1208 2813 -1184 2847
rect -1208 2779 -1162 2813
rect -1208 2745 -1184 2779
rect -1208 2711 -1162 2745
rect -1208 2677 -1184 2711
rect -1208 2643 -1162 2677
rect -1208 2609 -1184 2643
rect -1208 2575 -1162 2609
rect -1208 2541 -1184 2575
rect -1208 2507 -1162 2541
rect -1208 2473 -1184 2507
rect -1208 2439 -1162 2473
rect -1208 2405 -1184 2439
rect -1208 2371 -1162 2405
rect -1208 2337 -1184 2371
rect -1208 2303 -1162 2337
rect -1208 2269 -1184 2303
rect -1208 2235 -1162 2269
rect -1208 2201 -1184 2235
rect -1208 2167 -1162 2201
rect -1208 2133 -1184 2167
rect -1208 2099 -1162 2133
rect -1208 2065 -1184 2099
rect -1208 2031 -1162 2065
rect -1208 1997 -1184 2031
rect -1208 1963 -1162 1997
rect -1208 1929 -1184 1963
rect -1208 1895 -1162 1929
rect -1208 1861 -1184 1895
rect -1208 1827 -1162 1861
rect -1208 1793 -1184 1827
rect -1208 1759 -1162 1793
rect -1208 1725 -1184 1759
rect -1208 1691 -1162 1725
rect -1208 1657 -1184 1691
rect -1208 1623 -1162 1657
rect -1208 1589 -1184 1623
rect -1208 1555 -1162 1589
rect -1208 1521 -1184 1555
rect -1208 1487 -1162 1521
rect -1208 1453 -1184 1487
rect -1208 1419 -1162 1453
rect -1208 1385 -1184 1419
rect -1208 1351 -1162 1385
rect -1208 1317 -1184 1351
rect -1208 1283 -1162 1317
rect -1208 1249 -1184 1283
rect -1208 1215 -1162 1249
rect -1208 1181 -1184 1215
rect -1208 1147 -1162 1181
rect -1208 1113 -1184 1147
rect -1208 1079 -1162 1113
rect -1208 1045 -1184 1079
rect -1208 1011 -1162 1045
rect -1208 977 -1184 1011
rect -1208 943 -1162 977
rect -1208 909 -1184 943
rect -1208 875 -1162 909
rect -1208 841 -1184 875
rect -1208 807 -1162 841
rect -1208 773 -1184 807
rect -1208 739 -1162 773
rect -1208 705 -1184 739
rect -1208 671 -1162 705
rect -1208 637 -1184 671
rect -1208 603 -1162 637
rect -1208 569 -1184 603
rect -1208 535 -1162 569
rect -1208 501 -1184 535
rect -1208 467 -1162 501
rect -1208 433 -1184 467
rect -1208 399 -1162 433
rect -1208 365 -1184 399
rect -1208 331 -1162 365
rect -1208 297 -1184 331
rect -1208 263 -1162 297
rect -1208 229 -1184 263
rect -1208 195 -1162 229
rect -1208 161 -1184 195
rect -1208 127 -1162 161
rect -1208 93 -1184 127
rect -1208 59 -1162 93
rect -1208 25 -1184 59
rect -1208 -9 -1162 25
rect -1208 -43 -1184 -9
rect -1208 -77 -1162 -43
rect -1208 -111 -1184 -77
rect -1208 -145 -1162 -111
rect -1208 -179 -1184 -145
rect -1208 -213 -1162 -179
rect -1208 -247 -1184 -213
rect -1208 -281 -1162 -247
rect -1208 -315 -1184 -281
rect -1208 -349 -1162 -315
rect -1208 -383 -1184 -349
rect -1208 -417 -1162 -383
rect -1208 -451 -1184 -417
rect -1208 -485 -1162 -451
rect -1208 -519 -1184 -485
rect -1208 -553 -1162 -519
rect -1208 -587 -1184 -553
rect -1208 -621 -1162 -587
rect -1208 -655 -1184 -621
rect -1208 -689 -1162 -655
rect -1208 -723 -1184 -689
rect -1208 -757 -1162 -723
rect -1208 -791 -1184 -757
rect -1208 -825 -1162 -791
rect -1208 -859 -1184 -825
rect -1208 -893 -1162 -859
rect -1208 -927 -1184 -893
rect -912 -894 -896 6870
rect 0 5969 300 6000
rect 0 31 25 5969
rect 275 31 300 5969
rect 0 0 300 31
rect -189 -651 489 -649
rect -190 -665 489 -651
rect -190 -835 -173 -665
rect 473 -835 489 -665
rect -190 -894 489 -835
rect 1196 -894 1212 6870
rect 1462 6859 1508 6893
rect 1484 6825 1508 6859
rect 1462 6791 1508 6825
rect 1484 6757 1508 6791
rect 1462 6723 1508 6757
rect 1484 6689 1508 6723
rect 1462 6655 1508 6689
rect 1484 6621 1508 6655
rect 1462 6587 1508 6621
rect 1484 6553 1508 6587
rect 1462 6519 1508 6553
rect 1484 6485 1508 6519
rect 1462 6451 1508 6485
rect 1484 6417 1508 6451
rect 1462 6383 1508 6417
rect 1484 6349 1508 6383
rect 1462 6315 1508 6349
rect 1484 6281 1508 6315
rect 1462 6247 1508 6281
rect 1484 6213 1508 6247
rect 1462 6179 1508 6213
rect 1484 6145 1508 6179
rect 1462 6111 1508 6145
rect 1484 6077 1508 6111
rect 1462 6043 1508 6077
rect 1484 6009 1508 6043
rect 1462 5975 1508 6009
rect 1484 5941 1508 5975
rect 1462 5907 1508 5941
rect 1484 5873 1508 5907
rect 1462 5839 1508 5873
rect 1484 5805 1508 5839
rect 1462 5771 1508 5805
rect 1484 5737 1508 5771
rect 1462 5703 1508 5737
rect 1484 5669 1508 5703
rect 1462 5635 1508 5669
rect 1484 5601 1508 5635
rect 1462 5567 1508 5601
rect 1484 5533 1508 5567
rect 1462 5499 1508 5533
rect 1484 5465 1508 5499
rect 1462 5431 1508 5465
rect 1484 5397 1508 5431
rect 1462 5363 1508 5397
rect 1484 5329 1508 5363
rect 1462 5295 1508 5329
rect 1484 5261 1508 5295
rect 1462 5227 1508 5261
rect 1484 5193 1508 5227
rect 1462 5159 1508 5193
rect 1484 5125 1508 5159
rect 1462 5091 1508 5125
rect 1484 5057 1508 5091
rect 1462 5023 1508 5057
rect 1484 4989 1508 5023
rect 1462 4955 1508 4989
rect 1484 4921 1508 4955
rect 1462 4887 1508 4921
rect 1484 4853 1508 4887
rect 1462 4819 1508 4853
rect 1484 4785 1508 4819
rect 1462 4751 1508 4785
rect 1484 4717 1508 4751
rect 1462 4683 1508 4717
rect 1484 4649 1508 4683
rect 1462 4615 1508 4649
rect 1484 4581 1508 4615
rect 1462 4547 1508 4581
rect 1484 4513 1508 4547
rect 1462 4479 1508 4513
rect 1484 4445 1508 4479
rect 1462 4411 1508 4445
rect 1484 4377 1508 4411
rect 1462 4343 1508 4377
rect 1484 4309 1508 4343
rect 1462 4275 1508 4309
rect 1484 4241 1508 4275
rect 1462 4207 1508 4241
rect 1484 4173 1508 4207
rect 1462 4139 1508 4173
rect 1484 4105 1508 4139
rect 1462 4071 1508 4105
rect 1484 4037 1508 4071
rect 1462 4003 1508 4037
rect 1484 3969 1508 4003
rect 1462 3935 1508 3969
rect 1484 3901 1508 3935
rect 1462 3867 1508 3901
rect 1484 3833 1508 3867
rect 1462 3799 1508 3833
rect 1484 3765 1508 3799
rect 1462 3731 1508 3765
rect 1484 3697 1508 3731
rect 1462 3663 1508 3697
rect 1484 3629 1508 3663
rect 1462 3595 1508 3629
rect 1484 3561 1508 3595
rect 1462 3527 1508 3561
rect 1484 3493 1508 3527
rect 1462 3459 1508 3493
rect 1484 3425 1508 3459
rect 1462 3391 1508 3425
rect 1484 3357 1508 3391
rect 1462 3323 1508 3357
rect 1484 3289 1508 3323
rect 1462 3255 1508 3289
rect 1484 3221 1508 3255
rect 1462 3187 1508 3221
rect 1484 3153 1508 3187
rect 1462 3119 1508 3153
rect 1484 3085 1508 3119
rect 1462 3051 1508 3085
rect 1484 3017 1508 3051
rect 1462 2983 1508 3017
rect 1484 2949 1508 2983
rect 1462 2915 1508 2949
rect 1484 2881 1508 2915
rect 1462 2847 1508 2881
rect 1484 2813 1508 2847
rect 1462 2779 1508 2813
rect 1484 2745 1508 2779
rect 1462 2711 1508 2745
rect 1484 2677 1508 2711
rect 1462 2643 1508 2677
rect 1484 2609 1508 2643
rect 1462 2575 1508 2609
rect 1484 2541 1508 2575
rect 1462 2507 1508 2541
rect 1484 2473 1508 2507
rect 1462 2439 1508 2473
rect 1484 2405 1508 2439
rect 1462 2371 1508 2405
rect 1484 2337 1508 2371
rect 1462 2303 1508 2337
rect 1484 2269 1508 2303
rect 1462 2235 1508 2269
rect 1484 2201 1508 2235
rect 1462 2167 1508 2201
rect 1484 2133 1508 2167
rect 1462 2099 1508 2133
rect 1484 2065 1508 2099
rect 1462 2031 1508 2065
rect 1484 1997 1508 2031
rect 1462 1963 1508 1997
rect 1484 1929 1508 1963
rect 1462 1895 1508 1929
rect 1484 1861 1508 1895
rect 1462 1827 1508 1861
rect 1484 1793 1508 1827
rect 1462 1759 1508 1793
rect 1484 1725 1508 1759
rect 1462 1691 1508 1725
rect 1484 1657 1508 1691
rect 1462 1623 1508 1657
rect 1484 1589 1508 1623
rect 1462 1555 1508 1589
rect 1484 1521 1508 1555
rect 1462 1487 1508 1521
rect 1484 1453 1508 1487
rect 1462 1419 1508 1453
rect 1484 1385 1508 1419
rect 1462 1351 1508 1385
rect 1484 1317 1508 1351
rect 1462 1283 1508 1317
rect 1484 1249 1508 1283
rect 1462 1215 1508 1249
rect 1484 1181 1508 1215
rect 1462 1147 1508 1181
rect 1484 1113 1508 1147
rect 1462 1079 1508 1113
rect 1484 1045 1508 1079
rect 1462 1011 1508 1045
rect 1484 977 1508 1011
rect 1462 943 1508 977
rect 1484 909 1508 943
rect 1462 875 1508 909
rect 1484 841 1508 875
rect 1462 807 1508 841
rect 1484 773 1508 807
rect 1462 739 1508 773
rect 1484 705 1508 739
rect 1462 671 1508 705
rect 1484 637 1508 671
rect 1462 603 1508 637
rect 1484 569 1508 603
rect 1462 535 1508 569
rect 1484 501 1508 535
rect 1462 467 1508 501
rect 1484 433 1508 467
rect 1462 399 1508 433
rect 1484 365 1508 399
rect 1462 331 1508 365
rect 1484 297 1508 331
rect 1462 263 1508 297
rect 1484 229 1508 263
rect 1462 195 1508 229
rect 1484 161 1508 195
rect 1462 127 1508 161
rect 1484 93 1508 127
rect 1462 59 1508 93
rect 1484 25 1508 59
rect 1462 -9 1508 25
rect 1484 -43 1508 -9
rect 1462 -77 1508 -43
rect 1484 -111 1508 -77
rect 1462 -145 1508 -111
rect 1484 -179 1508 -145
rect 1462 -213 1508 -179
rect 1484 -247 1508 -213
rect 1462 -281 1508 -247
rect 1484 -315 1508 -281
rect 1462 -349 1508 -315
rect 1484 -383 1508 -349
rect 1462 -417 1508 -383
rect 1484 -451 1508 -417
rect 1462 -485 1508 -451
rect 1484 -519 1508 -485
rect 1462 -553 1508 -519
rect 1484 -587 1508 -553
rect 1462 -621 1508 -587
rect 1484 -655 1508 -621
rect 1462 -689 1508 -655
rect 1484 -723 1508 -689
rect 1462 -757 1508 -723
rect 1484 -791 1508 -757
rect 1462 -825 1508 -791
rect 1484 -859 1508 -825
rect 1462 -893 1508 -859
rect -912 -907 1212 -894
rect -1208 -961 -1162 -927
rect -1208 -995 -1184 -961
rect -1208 -1029 -1162 -995
rect -1208 -1063 -1184 -1029
rect -1208 -1157 -1162 -1063
rect -912 -1124 -839 -907
rect 1139 -1124 1212 -907
rect 1484 -927 1508 -893
rect 1462 -961 1508 -927
rect 1484 -995 1508 -961
rect 1462 -1029 1508 -995
rect 1484 -1063 1508 -1029
rect -912 -1157 -887 -1124
rect -1208 -1158 -1159 -1157
rect -1125 -1158 -1091 -1157
rect -1057 -1158 -1023 -1157
rect -989 -1158 -955 -1157
rect -921 -1158 -887 -1157
rect -853 -1157 -839 -1124
rect 1139 -1157 1153 -1124
rect -853 -1158 -819 -1157
rect -785 -1158 -751 -1157
rect -717 -1158 -683 -1157
rect -649 -1158 -615 -1157
rect -581 -1158 -547 -1157
rect -513 -1158 -479 -1157
rect -445 -1158 -411 -1157
rect -377 -1158 -343 -1157
rect -309 -1158 -275 -1157
rect -241 -1158 -207 -1157
rect -173 -1158 -139 -1157
rect -105 -1158 -71 -1157
rect -37 -1158 -3 -1157
rect 31 -1158 65 -1157
rect 99 -1158 133 -1157
rect 167 -1158 201 -1157
rect 235 -1158 269 -1157
rect 303 -1158 337 -1157
rect 371 -1158 405 -1157
rect 439 -1158 473 -1157
rect 507 -1158 541 -1157
rect 575 -1158 609 -1157
rect 643 -1158 677 -1157
rect 711 -1158 745 -1157
rect 779 -1158 813 -1157
rect 847 -1158 881 -1157
rect 915 -1158 949 -1157
rect 983 -1158 1017 -1157
rect 1051 -1158 1085 -1157
rect 1119 -1158 1153 -1157
rect 1187 -1157 1212 -1124
rect 1462 -1157 1508 -1063
rect 1187 -1158 1221 -1157
rect 1255 -1158 1289 -1157
rect 1323 -1158 1357 -1157
rect 1391 -1158 1425 -1157
rect 1459 -1158 1508 -1157
rect -1208 -1182 1508 -1158
<< viali >>
rect -1162 7124 -1159 7157
rect -1159 7124 -1125 7157
rect -1125 7124 -1091 7157
rect -1091 7124 -1057 7157
rect -1057 7124 -1023 7157
rect -1023 7124 -989 7157
rect -989 7124 -955 7157
rect -955 7124 -921 7157
rect -921 7124 -912 7157
rect -839 7124 -819 7157
rect -819 7124 -785 7157
rect -785 7124 -751 7157
rect -751 7124 -717 7157
rect -717 7124 -683 7157
rect -683 7124 -649 7157
rect -649 7124 -615 7157
rect -615 7124 -581 7157
rect -581 7124 -547 7157
rect -547 7124 -513 7157
rect -513 7124 -479 7157
rect -479 7124 -445 7157
rect -445 7124 -411 7157
rect -411 7124 -377 7157
rect -377 7124 -343 7157
rect -343 7124 -309 7157
rect -309 7124 -275 7157
rect -275 7124 -241 7157
rect -241 7124 -207 7157
rect -207 7124 -173 7157
rect -173 7124 -139 7157
rect -139 7124 -105 7157
rect -105 7124 -71 7157
rect -71 7124 -37 7157
rect -37 7124 -3 7157
rect -3 7124 31 7157
rect 31 7124 65 7157
rect 65 7124 99 7157
rect 99 7124 133 7157
rect 133 7124 167 7157
rect 167 7124 201 7157
rect 201 7124 235 7157
rect 235 7124 269 7157
rect 269 7124 303 7157
rect 303 7124 337 7157
rect 337 7124 371 7157
rect 371 7124 405 7157
rect 405 7124 439 7157
rect 439 7124 473 7157
rect 473 7124 507 7157
rect 507 7124 541 7157
rect 541 7124 575 7157
rect 575 7124 609 7157
rect 609 7124 643 7157
rect 643 7124 677 7157
rect 677 7124 711 7157
rect 711 7124 745 7157
rect 745 7124 779 7157
rect 779 7124 813 7157
rect 813 7124 847 7157
rect 847 7124 881 7157
rect 881 7124 915 7157
rect 915 7124 949 7157
rect 949 7124 983 7157
rect 983 7124 1017 7157
rect 1017 7124 1051 7157
rect 1051 7124 1085 7157
rect 1085 7124 1119 7157
rect 1119 7124 1139 7157
rect 1212 7124 1221 7157
rect 1221 7124 1255 7157
rect 1255 7124 1289 7157
rect 1289 7124 1323 7157
rect 1323 7124 1357 7157
rect 1357 7124 1391 7157
rect 1391 7124 1425 7157
rect 1425 7124 1459 7157
rect 1459 7124 1462 7157
rect -1162 7063 -912 7124
rect -1162 7029 -1150 7063
rect -1150 7029 -912 7063
rect -1162 6995 -912 7029
rect -1162 6961 -1150 6995
rect -1150 6961 -912 6995
rect -1162 6927 -912 6961
rect -1162 6893 -1150 6927
rect -1150 6893 -912 6927
rect -839 6907 1139 7124
rect 1212 7063 1462 7124
rect 1212 7029 1450 7063
rect 1450 7029 1462 7063
rect 1212 6995 1462 7029
rect 1212 6961 1450 6995
rect 1450 6961 1462 6995
rect 1212 6927 1462 6961
rect -1162 6859 -912 6893
rect 1212 6893 1450 6927
rect 1450 6893 1462 6927
rect -1162 6825 -1150 6859
rect -1150 6825 -912 6859
rect -1162 6791 -912 6825
rect -1162 6757 -1150 6791
rect -1150 6757 -912 6791
rect -1162 6723 -912 6757
rect -1162 6689 -1150 6723
rect -1150 6689 -912 6723
rect -1162 6655 -912 6689
rect -1162 6621 -1150 6655
rect -1150 6621 -912 6655
rect -1162 6587 -912 6621
rect -1162 6553 -1150 6587
rect -1150 6553 -912 6587
rect -1162 6519 -912 6553
rect -1162 6485 -1150 6519
rect -1150 6485 -912 6519
rect -1162 6451 -912 6485
rect -1162 6417 -1150 6451
rect -1150 6417 -912 6451
rect -1162 6383 -912 6417
rect -1162 6349 -1150 6383
rect -1150 6349 -912 6383
rect -1162 6315 -912 6349
rect -1162 6281 -1150 6315
rect -1150 6281 -912 6315
rect -1162 6247 -912 6281
rect -1162 6213 -1150 6247
rect -1150 6213 -912 6247
rect -1162 6179 -912 6213
rect -1162 6145 -1150 6179
rect -1150 6145 -912 6179
rect -1162 6111 -912 6145
rect -1162 6077 -1150 6111
rect -1150 6077 -912 6111
rect -1162 6043 -912 6077
rect -1162 6009 -1150 6043
rect -1150 6009 -912 6043
rect -1162 5975 -912 6009
rect -1162 5941 -1150 5975
rect -1150 5941 -1014 5975
rect -1162 5907 -1014 5941
rect -1162 5873 -1150 5907
rect -1150 5873 -1014 5907
rect -1162 5839 -1014 5873
rect -1162 5805 -1150 5839
rect -1150 5805 -1014 5839
rect -1162 5771 -1014 5805
rect -1162 5737 -1150 5771
rect -1150 5737 -1014 5771
rect -1162 5703 -1014 5737
rect -1162 5669 -1150 5703
rect -1150 5669 -1014 5703
rect -1162 5635 -1014 5669
rect -1162 5601 -1150 5635
rect -1150 5601 -1014 5635
rect -1162 5567 -1014 5601
rect -1162 5533 -1150 5567
rect -1150 5533 -1014 5567
rect -1162 5499 -1014 5533
rect -1162 5465 -1150 5499
rect -1150 5465 -1014 5499
rect -1162 5431 -1014 5465
rect -1162 5397 -1150 5431
rect -1150 5397 -1014 5431
rect -1162 5363 -1014 5397
rect -1162 5329 -1150 5363
rect -1150 5329 -1014 5363
rect -1162 5295 -1014 5329
rect -1162 5261 -1150 5295
rect -1150 5261 -1014 5295
rect -1162 5227 -1014 5261
rect -1162 5193 -1150 5227
rect -1150 5193 -1014 5227
rect -1162 5159 -1014 5193
rect -1162 5125 -1150 5159
rect -1150 5125 -1014 5159
rect -1162 5091 -1014 5125
rect -1162 5057 -1150 5091
rect -1150 5057 -1014 5091
rect -1162 5023 -1014 5057
rect -1162 4989 -1150 5023
rect -1150 4989 -1014 5023
rect -1162 4955 -1014 4989
rect -1162 4921 -1150 4955
rect -1150 4921 -1014 4955
rect -1162 4887 -1014 4921
rect -1162 4853 -1150 4887
rect -1150 4853 -1014 4887
rect -1162 4819 -1014 4853
rect -1162 4785 -1150 4819
rect -1150 4785 -1014 4819
rect -1162 4751 -1014 4785
rect -1162 4717 -1150 4751
rect -1150 4717 -1014 4751
rect -1162 4683 -1014 4717
rect -1162 4649 -1150 4683
rect -1150 4649 -1014 4683
rect -1162 4615 -1014 4649
rect -1162 4581 -1150 4615
rect -1150 4581 -1014 4615
rect -1162 4547 -1014 4581
rect -1162 4513 -1150 4547
rect -1150 4513 -1014 4547
rect -1162 4479 -1014 4513
rect -1162 4445 -1150 4479
rect -1150 4445 -1014 4479
rect -1162 4411 -1014 4445
rect -1162 4377 -1150 4411
rect -1150 4377 -1014 4411
rect -1162 4343 -1014 4377
rect -1162 4309 -1150 4343
rect -1150 4309 -1014 4343
rect -1162 4275 -1014 4309
rect -1162 4241 -1150 4275
rect -1150 4241 -1014 4275
rect -1162 4207 -1014 4241
rect -1162 4173 -1150 4207
rect -1150 4173 -1014 4207
rect -1162 4139 -1014 4173
rect -1162 4105 -1150 4139
rect -1150 4105 -1014 4139
rect -1162 4071 -1014 4105
rect -1162 4037 -1150 4071
rect -1150 4037 -1014 4071
rect -1162 4003 -1014 4037
rect -1162 3969 -1150 4003
rect -1150 3969 -1014 4003
rect -1162 3935 -1014 3969
rect -1162 3901 -1150 3935
rect -1150 3901 -1014 3935
rect -1162 3867 -1014 3901
rect -1162 3833 -1150 3867
rect -1150 3833 -1014 3867
rect -1162 3799 -1014 3833
rect -1162 3765 -1150 3799
rect -1150 3765 -1014 3799
rect -1162 3731 -1014 3765
rect -1162 3697 -1150 3731
rect -1150 3697 -1014 3731
rect -1162 3663 -1014 3697
rect -1162 3629 -1150 3663
rect -1150 3629 -1014 3663
rect -1162 3595 -1014 3629
rect -1162 3561 -1150 3595
rect -1150 3561 -1014 3595
rect -1162 3527 -1014 3561
rect -1162 3493 -1150 3527
rect -1150 3493 -1014 3527
rect -1162 3459 -1014 3493
rect -1162 3425 -1150 3459
rect -1150 3425 -1014 3459
rect -1162 3391 -1014 3425
rect -1162 3357 -1150 3391
rect -1150 3357 -1014 3391
rect -1162 3323 -1014 3357
rect -1162 3289 -1150 3323
rect -1150 3289 -1014 3323
rect -1162 3255 -1014 3289
rect -1162 3221 -1150 3255
rect -1150 3221 -1014 3255
rect -1162 3187 -1014 3221
rect -1162 3153 -1150 3187
rect -1150 3153 -1014 3187
rect -1162 3119 -1014 3153
rect -1162 3085 -1150 3119
rect -1150 3085 -1014 3119
rect -1162 3051 -1014 3085
rect -1162 3017 -1150 3051
rect -1150 3017 -1014 3051
rect -1162 2983 -1014 3017
rect -1162 2949 -1150 2983
rect -1150 2949 -1014 2983
rect -1162 2915 -1014 2949
rect -1162 2881 -1150 2915
rect -1150 2881 -1014 2915
rect -1162 2847 -1014 2881
rect -1162 2813 -1150 2847
rect -1150 2813 -1014 2847
rect -1162 2779 -1014 2813
rect -1162 2745 -1150 2779
rect -1150 2745 -1014 2779
rect -1162 2711 -1014 2745
rect -1162 2677 -1150 2711
rect -1150 2677 -1014 2711
rect -1162 2643 -1014 2677
rect -1162 2609 -1150 2643
rect -1150 2609 -1014 2643
rect -1162 2575 -1014 2609
rect -1162 2541 -1150 2575
rect -1150 2541 -1014 2575
rect -1162 2507 -1014 2541
rect -1162 2473 -1150 2507
rect -1150 2473 -1014 2507
rect -1162 2439 -1014 2473
rect -1162 2405 -1150 2439
rect -1150 2405 -1014 2439
rect -1162 2371 -1014 2405
rect -1162 2337 -1150 2371
rect -1150 2337 -1014 2371
rect -1162 2303 -1014 2337
rect -1162 2269 -1150 2303
rect -1150 2269 -1014 2303
rect -1162 2235 -1014 2269
rect -1162 2201 -1150 2235
rect -1150 2201 -1014 2235
rect -1162 2167 -1014 2201
rect -1162 2133 -1150 2167
rect -1150 2133 -1014 2167
rect -1162 2099 -1014 2133
rect -1162 2065 -1150 2099
rect -1150 2065 -1014 2099
rect -1162 2031 -1014 2065
rect -1162 1997 -1150 2031
rect -1150 1997 -1014 2031
rect -1162 1963 -1014 1997
rect -1162 1929 -1150 1963
rect -1150 1929 -1014 1963
rect -1162 1895 -1014 1929
rect -1162 1861 -1150 1895
rect -1150 1861 -1014 1895
rect -1162 1827 -1014 1861
rect -1162 1793 -1150 1827
rect -1150 1793 -1014 1827
rect -1162 1759 -1014 1793
rect -1162 1725 -1150 1759
rect -1150 1725 -1014 1759
rect -1162 1691 -1014 1725
rect -1162 1657 -1150 1691
rect -1150 1657 -1014 1691
rect -1162 1623 -1014 1657
rect -1162 1589 -1150 1623
rect -1150 1589 -1014 1623
rect -1162 1555 -1014 1589
rect -1162 1521 -1150 1555
rect -1150 1521 -1014 1555
rect -1162 1487 -1014 1521
rect -1162 1453 -1150 1487
rect -1150 1453 -1014 1487
rect -1162 1419 -1014 1453
rect -1162 1385 -1150 1419
rect -1150 1385 -1014 1419
rect -1162 1351 -1014 1385
rect -1162 1317 -1150 1351
rect -1150 1317 -1014 1351
rect -1162 1283 -1014 1317
rect -1162 1249 -1150 1283
rect -1150 1249 -1014 1283
rect -1162 1215 -1014 1249
rect -1162 1181 -1150 1215
rect -1150 1181 -1014 1215
rect -1162 1147 -1014 1181
rect -1162 1113 -1150 1147
rect -1150 1113 -1014 1147
rect -1162 1079 -1014 1113
rect -1162 1045 -1150 1079
rect -1150 1045 -1014 1079
rect -1162 1011 -1014 1045
rect -1162 977 -1150 1011
rect -1150 977 -1014 1011
rect -1162 943 -1014 977
rect -1162 909 -1150 943
rect -1150 909 -1014 943
rect -1162 875 -1014 909
rect -1162 841 -1150 875
rect -1150 841 -1014 875
rect -1162 807 -1014 841
rect -1162 773 -1150 807
rect -1150 773 -1014 807
rect -1162 739 -1014 773
rect -1162 705 -1150 739
rect -1150 705 -1014 739
rect -1162 671 -1014 705
rect -1162 637 -1150 671
rect -1150 637 -1014 671
rect -1162 603 -1014 637
rect -1162 569 -1150 603
rect -1150 569 -1014 603
rect -1162 535 -1014 569
rect -1162 501 -1150 535
rect -1150 501 -1014 535
rect -1162 467 -1014 501
rect -1162 433 -1150 467
rect -1150 433 -1014 467
rect -1162 399 -1014 433
rect -1162 365 -1150 399
rect -1150 365 -1014 399
rect -1162 331 -1014 365
rect -1162 297 -1150 331
rect -1150 297 -1014 331
rect -1162 263 -1014 297
rect -1162 229 -1150 263
rect -1150 229 -1014 263
rect -1162 195 -1014 229
rect -1162 161 -1150 195
rect -1150 161 -1014 195
rect -1162 127 -1014 161
rect -1162 93 -1150 127
rect -1150 93 -1014 127
rect -1162 59 -1014 93
rect -1162 25 -1150 59
rect -1150 25 -1014 59
rect -1014 25 -912 5975
rect -1162 -9 -912 25
rect -1162 -43 -1150 -9
rect -1150 -43 -912 -9
rect -1162 -77 -912 -43
rect -1162 -111 -1150 -77
rect -1150 -111 -912 -77
rect -1162 -145 -912 -111
rect -1162 -179 -1150 -145
rect -1150 -179 -912 -145
rect -1162 -213 -912 -179
rect -1162 -247 -1150 -213
rect -1150 -247 -912 -213
rect -1162 -281 -912 -247
rect -1162 -315 -1150 -281
rect -1150 -315 -912 -281
rect -1162 -349 -912 -315
rect -1162 -383 -1150 -349
rect -1150 -383 -912 -349
rect -1162 -417 -912 -383
rect -1162 -451 -1150 -417
rect -1150 -451 -912 -417
rect -1162 -485 -912 -451
rect -1162 -519 -1150 -485
rect -1150 -519 -912 -485
rect -1162 -553 -912 -519
rect -1162 -587 -1150 -553
rect -1150 -587 -912 -553
rect -1162 -621 -912 -587
rect -1162 -655 -1150 -621
rect -1150 -655 -912 -621
rect -1162 -689 -912 -655
rect -1162 -723 -1150 -689
rect -1150 -723 -912 -689
rect -1162 -757 -912 -723
rect -1162 -791 -1150 -757
rect -1150 -791 -912 -757
rect -1162 -825 -912 -791
rect -1162 -859 -1150 -825
rect -1150 -859 -912 -825
rect -1162 -893 -912 -859
rect -1162 -927 -1150 -893
rect -1150 -927 -912 -893
rect 25 5941 275 5969
rect 25 59 31 5941
rect 31 59 269 5941
rect 269 59 275 5941
rect 25 31 275 59
rect 1212 6859 1462 6893
rect 1212 6825 1450 6859
rect 1450 6825 1462 6859
rect 1212 6791 1462 6825
rect 1212 6757 1450 6791
rect 1450 6757 1462 6791
rect 1212 6723 1462 6757
rect 1212 6689 1450 6723
rect 1450 6689 1462 6723
rect 1212 6655 1462 6689
rect 1212 6621 1450 6655
rect 1450 6621 1462 6655
rect 1212 6587 1462 6621
rect 1212 6553 1450 6587
rect 1450 6553 1462 6587
rect 1212 6519 1462 6553
rect 1212 6485 1450 6519
rect 1450 6485 1462 6519
rect 1212 6451 1462 6485
rect 1212 6417 1450 6451
rect 1450 6417 1462 6451
rect 1212 6383 1462 6417
rect 1212 6349 1450 6383
rect 1450 6349 1462 6383
rect 1212 6315 1462 6349
rect 1212 6281 1450 6315
rect 1450 6281 1462 6315
rect 1212 6247 1462 6281
rect 1212 6213 1450 6247
rect 1450 6213 1462 6247
rect 1212 6179 1462 6213
rect 1212 6145 1450 6179
rect 1450 6145 1462 6179
rect 1212 6111 1462 6145
rect 1212 6077 1450 6111
rect 1450 6077 1462 6111
rect 1212 6043 1462 6077
rect 1212 6009 1450 6043
rect 1450 6009 1462 6043
rect 1212 5975 1462 6009
rect 1212 25 1314 5975
rect 1314 5941 1450 5975
rect 1450 5941 1462 5975
rect 1314 5907 1462 5941
rect 1314 5873 1450 5907
rect 1450 5873 1462 5907
rect 1314 5839 1462 5873
rect 1314 5805 1450 5839
rect 1450 5805 1462 5839
rect 1314 5771 1462 5805
rect 1314 5737 1450 5771
rect 1450 5737 1462 5771
rect 1314 5703 1462 5737
rect 1314 5669 1450 5703
rect 1450 5669 1462 5703
rect 1314 5635 1462 5669
rect 1314 5601 1450 5635
rect 1450 5601 1462 5635
rect 1314 5567 1462 5601
rect 1314 5533 1450 5567
rect 1450 5533 1462 5567
rect 1314 5499 1462 5533
rect 1314 5465 1450 5499
rect 1450 5465 1462 5499
rect 1314 5431 1462 5465
rect 1314 5397 1450 5431
rect 1450 5397 1462 5431
rect 1314 5363 1462 5397
rect 1314 5329 1450 5363
rect 1450 5329 1462 5363
rect 1314 5295 1462 5329
rect 1314 5261 1450 5295
rect 1450 5261 1462 5295
rect 1314 5227 1462 5261
rect 1314 5193 1450 5227
rect 1450 5193 1462 5227
rect 1314 5159 1462 5193
rect 1314 5125 1450 5159
rect 1450 5125 1462 5159
rect 1314 5091 1462 5125
rect 1314 5057 1450 5091
rect 1450 5057 1462 5091
rect 1314 5023 1462 5057
rect 1314 4989 1450 5023
rect 1450 4989 1462 5023
rect 1314 4955 1462 4989
rect 1314 4921 1450 4955
rect 1450 4921 1462 4955
rect 1314 4887 1462 4921
rect 1314 4853 1450 4887
rect 1450 4853 1462 4887
rect 1314 4819 1462 4853
rect 1314 4785 1450 4819
rect 1450 4785 1462 4819
rect 1314 4751 1462 4785
rect 1314 4717 1450 4751
rect 1450 4717 1462 4751
rect 1314 4683 1462 4717
rect 1314 4649 1450 4683
rect 1450 4649 1462 4683
rect 1314 4615 1462 4649
rect 1314 4581 1450 4615
rect 1450 4581 1462 4615
rect 1314 4547 1462 4581
rect 1314 4513 1450 4547
rect 1450 4513 1462 4547
rect 1314 4479 1462 4513
rect 1314 4445 1450 4479
rect 1450 4445 1462 4479
rect 1314 4411 1462 4445
rect 1314 4377 1450 4411
rect 1450 4377 1462 4411
rect 1314 4343 1462 4377
rect 1314 4309 1450 4343
rect 1450 4309 1462 4343
rect 1314 4275 1462 4309
rect 1314 4241 1450 4275
rect 1450 4241 1462 4275
rect 1314 4207 1462 4241
rect 1314 4173 1450 4207
rect 1450 4173 1462 4207
rect 1314 4139 1462 4173
rect 1314 4105 1450 4139
rect 1450 4105 1462 4139
rect 1314 4071 1462 4105
rect 1314 4037 1450 4071
rect 1450 4037 1462 4071
rect 1314 4003 1462 4037
rect 1314 3969 1450 4003
rect 1450 3969 1462 4003
rect 1314 3935 1462 3969
rect 1314 3901 1450 3935
rect 1450 3901 1462 3935
rect 1314 3867 1462 3901
rect 1314 3833 1450 3867
rect 1450 3833 1462 3867
rect 1314 3799 1462 3833
rect 1314 3765 1450 3799
rect 1450 3765 1462 3799
rect 1314 3731 1462 3765
rect 1314 3697 1450 3731
rect 1450 3697 1462 3731
rect 1314 3663 1462 3697
rect 1314 3629 1450 3663
rect 1450 3629 1462 3663
rect 1314 3595 1462 3629
rect 1314 3561 1450 3595
rect 1450 3561 1462 3595
rect 1314 3527 1462 3561
rect 1314 3493 1450 3527
rect 1450 3493 1462 3527
rect 1314 3459 1462 3493
rect 1314 3425 1450 3459
rect 1450 3425 1462 3459
rect 1314 3391 1462 3425
rect 1314 3357 1450 3391
rect 1450 3357 1462 3391
rect 1314 3323 1462 3357
rect 1314 3289 1450 3323
rect 1450 3289 1462 3323
rect 1314 3255 1462 3289
rect 1314 3221 1450 3255
rect 1450 3221 1462 3255
rect 1314 3187 1462 3221
rect 1314 3153 1450 3187
rect 1450 3153 1462 3187
rect 1314 3119 1462 3153
rect 1314 3085 1450 3119
rect 1450 3085 1462 3119
rect 1314 3051 1462 3085
rect 1314 3017 1450 3051
rect 1450 3017 1462 3051
rect 1314 2983 1462 3017
rect 1314 2949 1450 2983
rect 1450 2949 1462 2983
rect 1314 2915 1462 2949
rect 1314 2881 1450 2915
rect 1450 2881 1462 2915
rect 1314 2847 1462 2881
rect 1314 2813 1450 2847
rect 1450 2813 1462 2847
rect 1314 2779 1462 2813
rect 1314 2745 1450 2779
rect 1450 2745 1462 2779
rect 1314 2711 1462 2745
rect 1314 2677 1450 2711
rect 1450 2677 1462 2711
rect 1314 2643 1462 2677
rect 1314 2609 1450 2643
rect 1450 2609 1462 2643
rect 1314 2575 1462 2609
rect 1314 2541 1450 2575
rect 1450 2541 1462 2575
rect 1314 2507 1462 2541
rect 1314 2473 1450 2507
rect 1450 2473 1462 2507
rect 1314 2439 1462 2473
rect 1314 2405 1450 2439
rect 1450 2405 1462 2439
rect 1314 2371 1462 2405
rect 1314 2337 1450 2371
rect 1450 2337 1462 2371
rect 1314 2303 1462 2337
rect 1314 2269 1450 2303
rect 1450 2269 1462 2303
rect 1314 2235 1462 2269
rect 1314 2201 1450 2235
rect 1450 2201 1462 2235
rect 1314 2167 1462 2201
rect 1314 2133 1450 2167
rect 1450 2133 1462 2167
rect 1314 2099 1462 2133
rect 1314 2065 1450 2099
rect 1450 2065 1462 2099
rect 1314 2031 1462 2065
rect 1314 1997 1450 2031
rect 1450 1997 1462 2031
rect 1314 1963 1462 1997
rect 1314 1929 1450 1963
rect 1450 1929 1462 1963
rect 1314 1895 1462 1929
rect 1314 1861 1450 1895
rect 1450 1861 1462 1895
rect 1314 1827 1462 1861
rect 1314 1793 1450 1827
rect 1450 1793 1462 1827
rect 1314 1759 1462 1793
rect 1314 1725 1450 1759
rect 1450 1725 1462 1759
rect 1314 1691 1462 1725
rect 1314 1657 1450 1691
rect 1450 1657 1462 1691
rect 1314 1623 1462 1657
rect 1314 1589 1450 1623
rect 1450 1589 1462 1623
rect 1314 1555 1462 1589
rect 1314 1521 1450 1555
rect 1450 1521 1462 1555
rect 1314 1487 1462 1521
rect 1314 1453 1450 1487
rect 1450 1453 1462 1487
rect 1314 1419 1462 1453
rect 1314 1385 1450 1419
rect 1450 1385 1462 1419
rect 1314 1351 1462 1385
rect 1314 1317 1450 1351
rect 1450 1317 1462 1351
rect 1314 1283 1462 1317
rect 1314 1249 1450 1283
rect 1450 1249 1462 1283
rect 1314 1215 1462 1249
rect 1314 1181 1450 1215
rect 1450 1181 1462 1215
rect 1314 1147 1462 1181
rect 1314 1113 1450 1147
rect 1450 1113 1462 1147
rect 1314 1079 1462 1113
rect 1314 1045 1450 1079
rect 1450 1045 1462 1079
rect 1314 1011 1462 1045
rect 1314 977 1450 1011
rect 1450 977 1462 1011
rect 1314 943 1462 977
rect 1314 909 1450 943
rect 1450 909 1462 943
rect 1314 875 1462 909
rect 1314 841 1450 875
rect 1450 841 1462 875
rect 1314 807 1462 841
rect 1314 773 1450 807
rect 1450 773 1462 807
rect 1314 739 1462 773
rect 1314 705 1450 739
rect 1450 705 1462 739
rect 1314 671 1462 705
rect 1314 637 1450 671
rect 1450 637 1462 671
rect 1314 603 1462 637
rect 1314 569 1450 603
rect 1450 569 1462 603
rect 1314 535 1462 569
rect 1314 501 1450 535
rect 1450 501 1462 535
rect 1314 467 1462 501
rect 1314 433 1450 467
rect 1450 433 1462 467
rect 1314 399 1462 433
rect 1314 365 1450 399
rect 1450 365 1462 399
rect 1314 331 1462 365
rect 1314 297 1450 331
rect 1450 297 1462 331
rect 1314 263 1462 297
rect 1314 229 1450 263
rect 1450 229 1462 263
rect 1314 195 1462 229
rect 1314 161 1450 195
rect 1450 161 1462 195
rect 1314 127 1462 161
rect 1314 93 1450 127
rect 1450 93 1462 127
rect 1314 59 1462 93
rect 1314 25 1450 59
rect 1450 25 1462 59
rect 1212 -9 1462 25
rect 1212 -43 1450 -9
rect 1450 -43 1462 -9
rect 1212 -77 1462 -43
rect 1212 -111 1450 -77
rect 1450 -111 1462 -77
rect 1212 -145 1462 -111
rect 1212 -179 1450 -145
rect 1450 -179 1462 -145
rect 1212 -213 1462 -179
rect 1212 -247 1450 -213
rect 1450 -247 1462 -213
rect 1212 -281 1462 -247
rect 1212 -315 1450 -281
rect 1450 -315 1462 -281
rect 1212 -349 1462 -315
rect 1212 -383 1450 -349
rect 1450 -383 1462 -349
rect 1212 -417 1462 -383
rect 1212 -451 1450 -417
rect 1450 -451 1462 -417
rect 1212 -485 1462 -451
rect 1212 -519 1450 -485
rect 1450 -519 1462 -485
rect 1212 -553 1462 -519
rect 1212 -587 1450 -553
rect 1450 -587 1462 -553
rect 1212 -621 1462 -587
rect 1212 -655 1450 -621
rect 1450 -655 1462 -621
rect 1212 -689 1462 -655
rect 1212 -723 1450 -689
rect 1450 -723 1462 -689
rect 1212 -757 1462 -723
rect 1212 -791 1450 -757
rect 1450 -791 1462 -757
rect 1212 -825 1462 -791
rect 1212 -859 1450 -825
rect 1450 -859 1462 -825
rect 1212 -893 1462 -859
rect -1162 -961 -912 -927
rect -1162 -995 -1150 -961
rect -1150 -995 -912 -961
rect -1162 -1029 -912 -995
rect -1162 -1063 -1150 -1029
rect -1150 -1063 -912 -1029
rect -1162 -1124 -912 -1063
rect -839 -1124 1139 -907
rect 1212 -927 1450 -893
rect 1450 -927 1462 -893
rect 1212 -961 1462 -927
rect 1212 -995 1450 -961
rect 1450 -995 1462 -961
rect 1212 -1029 1462 -995
rect 1212 -1063 1450 -1029
rect 1450 -1063 1462 -1029
rect 1212 -1124 1462 -1063
rect -1162 -1157 -1159 -1124
rect -1159 -1157 -1125 -1124
rect -1125 -1157 -1091 -1124
rect -1091 -1157 -1057 -1124
rect -1057 -1157 -1023 -1124
rect -1023 -1157 -989 -1124
rect -989 -1157 -955 -1124
rect -955 -1157 -921 -1124
rect -921 -1157 -912 -1124
rect -839 -1157 -819 -1124
rect -819 -1157 -785 -1124
rect -785 -1157 -751 -1124
rect -751 -1157 -717 -1124
rect -717 -1157 -683 -1124
rect -683 -1157 -649 -1124
rect -649 -1157 -615 -1124
rect -615 -1157 -581 -1124
rect -581 -1157 -547 -1124
rect -547 -1157 -513 -1124
rect -513 -1157 -479 -1124
rect -479 -1157 -445 -1124
rect -445 -1157 -411 -1124
rect -411 -1157 -377 -1124
rect -377 -1157 -343 -1124
rect -343 -1157 -309 -1124
rect -309 -1157 -275 -1124
rect -275 -1157 -241 -1124
rect -241 -1157 -207 -1124
rect -207 -1157 -173 -1124
rect -173 -1157 -139 -1124
rect -139 -1157 -105 -1124
rect -105 -1157 -71 -1124
rect -71 -1157 -37 -1124
rect -37 -1157 -3 -1124
rect -3 -1157 31 -1124
rect 31 -1157 65 -1124
rect 65 -1157 99 -1124
rect 99 -1157 133 -1124
rect 133 -1157 167 -1124
rect 167 -1157 201 -1124
rect 201 -1157 235 -1124
rect 235 -1157 269 -1124
rect 269 -1157 303 -1124
rect 303 -1157 337 -1124
rect 337 -1157 371 -1124
rect 371 -1157 405 -1124
rect 405 -1157 439 -1124
rect 439 -1157 473 -1124
rect 473 -1157 507 -1124
rect 507 -1157 541 -1124
rect 541 -1157 575 -1124
rect 575 -1157 609 -1124
rect 609 -1157 643 -1124
rect 643 -1157 677 -1124
rect 677 -1157 711 -1124
rect 711 -1157 745 -1124
rect 745 -1157 779 -1124
rect 779 -1157 813 -1124
rect 813 -1157 847 -1124
rect 847 -1157 881 -1124
rect 881 -1157 915 -1124
rect 915 -1157 949 -1124
rect 949 -1157 983 -1124
rect 983 -1157 1017 -1124
rect 1017 -1157 1051 -1124
rect 1051 -1157 1085 -1124
rect 1085 -1157 1119 -1124
rect 1119 -1157 1139 -1124
rect 1212 -1157 1221 -1124
rect 1221 -1157 1255 -1124
rect 1255 -1157 1289 -1124
rect 1289 -1157 1323 -1124
rect 1323 -1157 1357 -1124
rect 1357 -1157 1391 -1124
rect 1391 -1157 1425 -1124
rect 1425 -1157 1459 -1124
rect 1459 -1157 1462 -1124
<< metal1 >>
rect -1208 7157 1508 7182
rect -1208 7156 -1162 7157
rect -912 7156 -839 7157
rect 1139 7156 1212 7157
rect 1462 7156 1508 7157
rect -1208 -1152 -1186 7156
rect -750 6720 -708 6907
rect 1008 6720 1050 6907
rect -750 6700 1050 6720
rect -750 6450 -607 6700
tri -607 6450 -357 6700 nw
tri 658 6450 908 6700 ne
rect 908 6450 1050 6700
rect -750 -374 -709 6450
tri -709 6348 -607 6450 nw
tri -431 6392 -373 6450 se
rect -373 6392 674 6450
tri 674 6392 732 6450 sw
tri 908 6392 966 6450 ne
rect 966 6392 1050 6450
tri -449 6374 -431 6392 se
rect -431 6386 732 6392
rect -431 6374 -388 6386
tri -709 -374 -683 -348 sw
rect -449 -374 -388 6374
rect 688 6374 732 6386
tri 732 6374 750 6392 sw
rect -750 -450 -683 -374
tri -683 -450 -607 -374 sw
tri -449 -392 -431 -374 ne
rect -431 -386 -388 -374
rect 688 -374 750 6374
tri 966 6348 1010 6392 ne
tri 984 -374 1010 -348 se
rect 1010 -374 1050 6392
rect 688 -386 732 -374
rect -431 -392 732 -386
tri 732 -392 750 -374 nw
tri 966 -392 984 -374 se
rect 984 -392 1050 -374
tri -431 -450 -373 -392 ne
rect -373 -450 674 -392
tri 674 -450 732 -392 nw
tri 908 -450 966 -392 se
rect 966 -450 1050 -392
rect -750 -700 -607 -450
tri -607 -700 -357 -450 sw
tri 658 -700 908 -450 se
rect 908 -700 1050 -450
rect -750 -716 1050 -700
rect -750 -907 -708 -716
rect 1008 -907 1050 -716
rect 1486 -1152 1508 7156
rect -1208 -1157 -1162 -1152
rect -912 -1157 -839 -1152
rect 1139 -1157 1212 -1152
rect 1462 -1157 1508 -1152
rect -1208 -1182 1508 -1157
<< via1 >>
rect -1186 -1152 -1162 7156
rect -1162 -1152 -912 7156
rect -912 6907 -839 7156
rect -839 6907 -750 7156
rect -708 6907 1008 7156
rect 1050 6907 1139 7156
rect 1139 6907 1212 7156
rect -912 -907 -750 6907
rect -708 6720 1008 6907
rect -388 5969 688 6386
rect -388 31 25 5969
rect 25 31 275 5969
rect 275 31 688 5969
rect -388 -386 688 31
rect -708 -907 1008 -716
rect 1050 -907 1212 6907
rect -912 -1152 -839 -907
rect -839 -1152 -750 -907
rect -708 -1152 1008 -907
rect 1050 -1152 1139 -907
rect 1139 -1152 1212 -907
rect 1212 -1152 1462 7156
rect 1462 -1152 1486 7156
<< metal2 >>
rect -1208 7156 1508 7182
rect -1208 -1152 -1186 7156
rect -750 6720 -708 7156
rect 1008 6720 1050 7156
rect -750 6700 1050 6720
rect -750 6450 -607 6700
tri -607 6450 -357 6700 nw
tri 658 6450 908 6700 ne
rect 908 6450 1050 6700
rect -750 6386 -671 6450
tri -671 6386 -607 6450 nw
tri -426 6397 -373 6450 se
rect -373 6397 674 6450
tri 674 6397 727 6450 sw
tri 908 6397 961 6450 ne
rect 961 6397 1050 6450
tri -437 6386 -426 6397 se
rect -426 6388 727 6397
rect -426 6386 -397 6388
rect -750 -386 -709 6386
tri -709 6348 -671 6386 nw
tri -449 6374 -437 6386 se
rect -437 6374 -397 6386
tri -709 -386 -671 -348 sw
rect -449 -374 -397 6374
tri -449 -386 -437 -374 ne
rect -437 -386 -397 -374
rect 699 6374 727 6388
tri 727 6374 750 6397 sw
rect 699 -374 750 6374
tri 961 6348 1010 6397 ne
rect -750 -450 -671 -386
tri -671 -450 -607 -386 sw
tri -437 -397 -426 -386 ne
rect -426 -388 -397 -386
rect 699 -388 727 -374
rect -426 -397 727 -388
tri 727 -397 750 -374 nw
tri 961 -397 1010 -348 se
rect 1010 -397 1050 6397
tri -426 -450 -373 -397 ne
rect -373 -450 674 -397
tri 674 -450 727 -397 nw
tri 908 -450 961 -397 se
rect 961 -450 1050 -397
rect -750 -700 -607 -450
tri -607 -700 -357 -450 sw
tri 658 -700 908 -450 se
rect 908 -700 1050 -450
rect -750 -716 1050 -700
rect -750 -1152 -708 -716
rect 1008 -1152 1050 -716
rect 1486 -1152 1508 7156
rect -1208 -1182 1508 -1152
<< via2 >>
rect -397 6386 699 6388
rect -397 -386 -388 6386
rect -388 -386 688 6386
rect 688 -386 699 6386
rect -397 -388 699 -386
<< metal3 >>
rect -1208 6388 1508 7182
rect -1208 5182 -397 6388
rect -968 818 -397 5182
rect -1208 -388 -397 818
rect 699 5182 1508 6388
rect 699 818 1268 5182
rect 699 -388 1508 818
rect -1208 -1182 1508 -388
<< properties >>
string GDS_END 4415914
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3915686
<< end >>
