magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect 3770 6536 6467 7237
rect 3805 5999 6467 6536
rect 3900 5111 5249 5153
rect 3900 4350 6467 5111
rect 3867 3857 6467 4350
rect 3867 3750 5105 3857
rect -9346 2317 -8425 3018
<< pwell >>
rect 3845 7556 6259 7642
rect 3845 7342 6255 7556
rect 3842 5680 6255 5894
rect 3842 5594 6280 5680
rect 3940 5323 5098 5594
rect 5298 5447 6280 5594
rect 5314 5216 6244 5447
rect 3907 3538 5065 3580
rect 5286 3538 6271 3752
rect 3907 3452 6291 3538
rect 3907 3388 5174 3452
rect 5088 3358 5174 3388
rect -9309 2020 -8500 2212
<< mvnmos >>
rect 3924 7368 4044 7508
rect 4100 7368 4220 7508
rect 4400 7368 4520 7508
rect 4576 7368 4696 7508
rect 4752 7368 4872 7508
rect 4928 7368 5048 7508
rect 5228 7368 5348 7508
rect 5404 7368 5524 7508
rect 5704 7368 5824 7508
rect 5880 7368 6000 7508
rect 6056 7368 6176 7508
rect 3924 5728 4044 5868
rect 4100 5728 4220 5868
rect 4400 5728 4520 5868
rect 4576 5728 4696 5868
rect 4876 5728 4996 5868
rect 5052 5728 5172 5868
rect 5228 5728 5348 5868
rect 5404 5728 5524 5868
rect 5704 5728 5824 5868
rect 5880 5728 6000 5868
rect 6056 5728 6176 5868
rect 4019 5349 4139 5489
rect 4195 5349 4315 5489
rect 4371 5349 4491 5489
rect 4547 5349 4667 5489
rect 4723 5349 4843 5489
rect 4899 5349 5019 5489
rect 5393 5242 5513 5382
rect 5693 5242 5813 5382
rect 5869 5242 5989 5382
rect 6045 5242 6165 5382
rect 5368 3586 5488 3726
rect 5544 3586 5664 3726
rect 5720 3586 5840 3726
rect 5896 3586 6016 3726
rect 6072 3586 6192 3726
rect 3986 3414 4106 3554
rect 4162 3414 4282 3554
rect 4338 3414 4458 3554
rect 4514 3414 4634 3554
rect 4690 3414 4810 3554
rect 4866 3414 4986 3554
rect -9227 2046 -9107 2186
rect -9051 2046 -8931 2186
rect -8875 2046 -8755 2186
rect -8699 2046 -8579 2186
<< mvpmos >>
rect 3924 6970 4044 7170
rect 4100 6970 4220 7170
rect 4400 6970 4520 7170
rect 4576 6970 4696 7170
rect 4752 6970 4872 7170
rect 4928 6970 5048 7170
rect 5228 6970 5348 7170
rect 5404 6970 5524 7170
rect 5704 6970 5824 7170
rect 5880 6970 6000 7170
rect 6056 6970 6176 7170
rect 3924 6702 4044 6902
rect 4100 6702 4220 6902
rect 4400 6702 4520 6902
rect 4576 6702 4696 6902
rect 4752 6702 4872 6902
rect 4928 6702 5048 6902
rect 5228 6702 5348 6902
rect 5404 6702 5524 6902
rect 5704 6702 5824 6902
rect 5880 6702 6000 6902
rect 6056 6702 6176 6902
rect 3924 6334 4044 6534
rect 4100 6334 4220 6534
rect 4400 6334 4520 6534
rect 4576 6334 4696 6534
rect 4876 6334 4996 6534
rect 5052 6334 5172 6534
rect 5228 6334 5348 6534
rect 5404 6334 5524 6534
rect 5704 6334 5824 6534
rect 5880 6334 6000 6534
rect 6056 6334 6176 6534
rect 3924 6066 4044 6266
rect 4100 6066 4220 6266
rect 4400 6066 4520 6266
rect 4576 6066 4696 6266
rect 4876 6066 4996 6266
rect 5052 6066 5172 6266
rect 5228 6066 5348 6266
rect 5404 6066 5524 6266
rect 5704 6066 5824 6266
rect 5880 6066 6000 6266
rect 6056 6066 6176 6266
rect 4019 4887 4139 5087
rect 4195 4887 4315 5087
rect 4371 4887 4491 5087
rect 4547 4887 4667 5087
rect 4723 4887 4843 5087
rect 4899 4887 5019 5087
rect 5393 4844 5513 5044
rect 5693 4844 5813 5044
rect 5869 4844 5989 5044
rect 6045 4844 6165 5044
rect 4019 4619 4139 4819
rect 4195 4619 4315 4819
rect 4371 4619 4491 4819
rect 4547 4619 4667 4819
rect 4723 4619 4843 4819
rect 4899 4619 5019 4819
rect 5393 4576 5513 4776
rect 5693 4576 5813 4776
rect 5869 4576 5989 4776
rect 6045 4576 6165 4776
rect 3986 4084 4106 4284
rect 4162 4084 4282 4284
rect 4338 4084 4458 4284
rect 4514 4084 4634 4284
rect 4690 4084 4810 4284
rect 4866 4084 4986 4284
rect 5368 4192 5488 4392
rect 5544 4192 5664 4392
rect 5720 4192 5840 4392
rect 5896 4192 6016 4392
rect 6072 4192 6192 4392
rect 3986 3816 4106 4016
rect 4162 3816 4282 4016
rect 4338 3816 4458 4016
rect 4514 3816 4634 4016
rect 4690 3816 4810 4016
rect 4866 3816 4986 4016
rect 5368 3924 5488 4124
rect 5544 3924 5664 4124
rect 5720 3924 5840 4124
rect 5896 3924 6016 4124
rect 6072 3924 6192 4124
rect -9227 2652 -9107 2852
rect -9051 2652 -8931 2852
rect -8875 2652 -8755 2852
rect -8699 2652 -8579 2852
rect -9227 2384 -9107 2584
rect -9051 2384 -8931 2584
rect -8875 2384 -8755 2584
rect -8699 2384 -8579 2584
<< mvndiff >>
rect 3871 7482 3924 7508
rect 3871 7448 3879 7482
rect 3913 7448 3924 7482
rect 3871 7414 3924 7448
rect 3871 7380 3879 7414
rect 3913 7380 3924 7414
rect 3871 7368 3924 7380
rect 4044 7368 4100 7508
rect 4220 7482 4273 7508
rect 4220 7448 4231 7482
rect 4265 7448 4273 7482
rect 4220 7414 4273 7448
rect 4220 7380 4231 7414
rect 4265 7380 4273 7414
rect 4220 7368 4273 7380
rect 4347 7482 4400 7508
rect 4347 7448 4355 7482
rect 4389 7448 4400 7482
rect 4347 7414 4400 7448
rect 4347 7380 4355 7414
rect 4389 7380 4400 7414
rect 4347 7368 4400 7380
rect 4520 7368 4576 7508
rect 4696 7482 4752 7508
rect 4696 7448 4707 7482
rect 4741 7448 4752 7482
rect 4696 7414 4752 7448
rect 4696 7380 4707 7414
rect 4741 7380 4752 7414
rect 4696 7368 4752 7380
rect 4872 7368 4928 7508
rect 5048 7482 5101 7508
rect 5048 7448 5059 7482
rect 5093 7448 5101 7482
rect 5048 7414 5101 7448
rect 5048 7380 5059 7414
rect 5093 7380 5101 7414
rect 5048 7368 5101 7380
rect 5175 7482 5228 7508
rect 5175 7448 5183 7482
rect 5217 7448 5228 7482
rect 5175 7414 5228 7448
rect 5175 7380 5183 7414
rect 5217 7380 5228 7414
rect 5175 7368 5228 7380
rect 5348 7368 5404 7508
rect 5524 7482 5577 7508
rect 5524 7448 5535 7482
rect 5569 7448 5577 7482
rect 5524 7414 5577 7448
rect 5524 7380 5535 7414
rect 5569 7380 5577 7414
rect 5524 7368 5577 7380
rect 5651 7482 5704 7508
rect 5651 7448 5659 7482
rect 5693 7448 5704 7482
rect 5651 7414 5704 7448
rect 5651 7380 5659 7414
rect 5693 7380 5704 7414
rect 5651 7368 5704 7380
rect 5824 7482 5880 7508
rect 5824 7448 5835 7482
rect 5869 7448 5880 7482
rect 5824 7414 5880 7448
rect 5824 7380 5835 7414
rect 5869 7380 5880 7414
rect 5824 7368 5880 7380
rect 6000 7482 6056 7508
rect 6000 7448 6011 7482
rect 6045 7448 6056 7482
rect 6000 7414 6056 7448
rect 6000 7380 6011 7414
rect 6045 7380 6056 7414
rect 6000 7368 6056 7380
rect 6176 7482 6229 7508
rect 6176 7448 6187 7482
rect 6221 7448 6229 7482
rect 6176 7414 6229 7448
rect 6176 7380 6187 7414
rect 6221 7380 6229 7414
rect 6176 7368 6229 7380
rect 3868 5856 3924 5868
rect 3868 5822 3879 5856
rect 3913 5822 3924 5856
rect 3868 5788 3924 5822
rect 3868 5754 3879 5788
rect 3913 5754 3924 5788
rect 3868 5728 3924 5754
rect 4044 5856 4100 5868
rect 4044 5822 4055 5856
rect 4089 5822 4100 5856
rect 4044 5788 4100 5822
rect 4044 5754 4055 5788
rect 4089 5754 4100 5788
rect 4044 5728 4100 5754
rect 4220 5856 4273 5868
rect 4220 5822 4231 5856
rect 4265 5822 4273 5856
rect 4220 5788 4273 5822
rect 4220 5754 4231 5788
rect 4265 5754 4273 5788
rect 4220 5728 4273 5754
rect 4347 5856 4400 5868
rect 4347 5822 4355 5856
rect 4389 5822 4400 5856
rect 4347 5788 4400 5822
rect 4347 5754 4355 5788
rect 4389 5754 4400 5788
rect 4347 5728 4400 5754
rect 4520 5728 4576 5868
rect 4696 5856 4749 5868
rect 4696 5822 4707 5856
rect 4741 5822 4749 5856
rect 4696 5788 4749 5822
rect 4696 5754 4707 5788
rect 4741 5754 4749 5788
rect 4696 5728 4749 5754
rect 4823 5856 4876 5868
rect 4823 5822 4831 5856
rect 4865 5822 4876 5856
rect 4823 5788 4876 5822
rect 4823 5754 4831 5788
rect 4865 5754 4876 5788
rect 4823 5728 4876 5754
rect 4996 5728 5052 5868
rect 5172 5856 5228 5868
rect 5172 5822 5183 5856
rect 5217 5822 5228 5856
rect 5172 5788 5228 5822
rect 5172 5754 5183 5788
rect 5217 5754 5228 5788
rect 5172 5728 5228 5754
rect 5348 5728 5404 5868
rect 5524 5856 5577 5868
rect 5524 5822 5535 5856
rect 5569 5822 5577 5856
rect 5524 5788 5577 5822
rect 5524 5754 5535 5788
rect 5569 5754 5577 5788
rect 5524 5728 5577 5754
rect 5651 5856 5704 5868
rect 5651 5822 5659 5856
rect 5693 5822 5704 5856
rect 5651 5788 5704 5822
rect 5651 5754 5659 5788
rect 5693 5754 5704 5788
rect 5651 5728 5704 5754
rect 5824 5856 5880 5868
rect 5824 5822 5835 5856
rect 5869 5822 5880 5856
rect 5824 5788 5880 5822
rect 5824 5754 5835 5788
rect 5869 5754 5880 5788
rect 5824 5728 5880 5754
rect 6000 5856 6056 5868
rect 6000 5822 6011 5856
rect 6045 5822 6056 5856
rect 6000 5788 6056 5822
rect 6000 5754 6011 5788
rect 6045 5754 6056 5788
rect 6000 5728 6056 5754
rect 6176 5856 6229 5868
rect 6176 5822 6187 5856
rect 6221 5822 6229 5856
rect 6176 5788 6229 5822
rect 6176 5754 6187 5788
rect 6221 5754 6229 5788
rect 6176 5728 6229 5754
rect 3966 5477 4019 5489
rect 3966 5443 3974 5477
rect 4008 5443 4019 5477
rect 3966 5409 4019 5443
rect 3966 5375 3974 5409
rect 4008 5375 4019 5409
rect 3966 5349 4019 5375
rect 4139 5477 4195 5489
rect 4139 5443 4150 5477
rect 4184 5443 4195 5477
rect 4139 5409 4195 5443
rect 4139 5375 4150 5409
rect 4184 5375 4195 5409
rect 4139 5349 4195 5375
rect 4315 5477 4371 5489
rect 4315 5443 4326 5477
rect 4360 5443 4371 5477
rect 4315 5409 4371 5443
rect 4315 5375 4326 5409
rect 4360 5375 4371 5409
rect 4315 5349 4371 5375
rect 4491 5477 4547 5489
rect 4491 5443 4502 5477
rect 4536 5443 4547 5477
rect 4491 5409 4547 5443
rect 4491 5375 4502 5409
rect 4536 5375 4547 5409
rect 4491 5349 4547 5375
rect 4667 5477 4723 5489
rect 4667 5443 4678 5477
rect 4712 5443 4723 5477
rect 4667 5409 4723 5443
rect 4667 5375 4678 5409
rect 4712 5375 4723 5409
rect 4667 5349 4723 5375
rect 4843 5477 4899 5489
rect 4843 5443 4854 5477
rect 4888 5443 4899 5477
rect 4843 5409 4899 5443
rect 4843 5375 4854 5409
rect 4888 5375 4899 5409
rect 4843 5349 4899 5375
rect 5019 5477 5072 5489
rect 5019 5443 5030 5477
rect 5064 5443 5072 5477
rect 5019 5409 5072 5443
rect 5019 5375 5030 5409
rect 5064 5375 5072 5409
rect 5019 5349 5072 5375
rect 5340 5356 5393 5382
rect 5340 5322 5348 5356
rect 5382 5322 5393 5356
rect 5340 5288 5393 5322
rect 5340 5254 5348 5288
rect 5382 5254 5393 5288
rect 5340 5242 5393 5254
rect 5513 5356 5566 5382
rect 5513 5322 5524 5356
rect 5558 5322 5566 5356
rect 5513 5288 5566 5322
rect 5513 5254 5524 5288
rect 5558 5254 5566 5288
rect 5513 5242 5566 5254
rect 5640 5356 5693 5382
rect 5640 5322 5648 5356
rect 5682 5322 5693 5356
rect 5640 5288 5693 5322
rect 5640 5254 5648 5288
rect 5682 5254 5693 5288
rect 5640 5242 5693 5254
rect 5813 5356 5869 5382
rect 5813 5322 5824 5356
rect 5858 5322 5869 5356
rect 5813 5288 5869 5322
rect 5813 5254 5824 5288
rect 5858 5254 5869 5288
rect 5813 5242 5869 5254
rect 5989 5356 6045 5382
rect 5989 5322 6000 5356
rect 6034 5322 6045 5356
rect 5989 5288 6045 5322
rect 5989 5254 6000 5288
rect 6034 5254 6045 5288
rect 5989 5242 6045 5254
rect 6165 5356 6218 5382
rect 6165 5322 6176 5356
rect 6210 5322 6218 5356
rect 6165 5288 6218 5322
rect 6165 5254 6176 5288
rect 6210 5254 6218 5288
rect 6165 5242 6218 5254
rect 5312 3714 5368 3726
rect 5312 3680 5323 3714
rect 5357 3680 5368 3714
rect 5312 3646 5368 3680
rect 5312 3612 5323 3646
rect 5357 3612 5368 3646
rect 5312 3586 5368 3612
rect 5488 3714 5544 3726
rect 5488 3680 5499 3714
rect 5533 3680 5544 3714
rect 5488 3646 5544 3680
rect 5488 3612 5499 3646
rect 5533 3612 5544 3646
rect 5488 3586 5544 3612
rect 5664 3714 5720 3726
rect 5664 3680 5675 3714
rect 5709 3680 5720 3714
rect 5664 3646 5720 3680
rect 5664 3612 5675 3646
rect 5709 3612 5720 3646
rect 5664 3586 5720 3612
rect 5840 3714 5896 3726
rect 5840 3680 5851 3714
rect 5885 3680 5896 3714
rect 5840 3646 5896 3680
rect 5840 3612 5851 3646
rect 5885 3612 5896 3646
rect 5840 3586 5896 3612
rect 6016 3714 6072 3726
rect 6016 3680 6027 3714
rect 6061 3680 6072 3714
rect 6016 3646 6072 3680
rect 6016 3612 6027 3646
rect 6061 3612 6072 3646
rect 6016 3586 6072 3612
rect 6192 3714 6245 3726
rect 6192 3680 6203 3714
rect 6237 3680 6245 3714
rect 6192 3646 6245 3680
rect 6192 3612 6203 3646
rect 6237 3612 6245 3646
rect 6192 3586 6245 3612
rect 3933 3528 3986 3554
rect 3933 3494 3941 3528
rect 3975 3494 3986 3528
rect 3933 3460 3986 3494
rect 3933 3426 3941 3460
rect 3975 3426 3986 3460
rect 3933 3414 3986 3426
rect 4106 3528 4162 3554
rect 4106 3494 4117 3528
rect 4151 3494 4162 3528
rect 4106 3460 4162 3494
rect 4106 3426 4117 3460
rect 4151 3426 4162 3460
rect 4106 3414 4162 3426
rect 4282 3528 4338 3554
rect 4282 3494 4293 3528
rect 4327 3494 4338 3528
rect 4282 3460 4338 3494
rect 4282 3426 4293 3460
rect 4327 3426 4338 3460
rect 4282 3414 4338 3426
rect 4458 3528 4514 3554
rect 4458 3494 4469 3528
rect 4503 3494 4514 3528
rect 4458 3460 4514 3494
rect 4458 3426 4469 3460
rect 4503 3426 4514 3460
rect 4458 3414 4514 3426
rect 4634 3528 4690 3554
rect 4634 3494 4645 3528
rect 4679 3494 4690 3528
rect 4634 3460 4690 3494
rect 4634 3426 4645 3460
rect 4679 3426 4690 3460
rect 4634 3414 4690 3426
rect 4810 3528 4866 3554
rect 4810 3494 4821 3528
rect 4855 3494 4866 3528
rect 4810 3460 4866 3494
rect 4810 3426 4821 3460
rect 4855 3426 4866 3460
rect 4810 3414 4866 3426
rect 4986 3528 5039 3554
rect 4986 3494 4997 3528
rect 5031 3494 5039 3528
rect 4986 3460 5039 3494
rect 4986 3426 4997 3460
rect 5031 3426 5039 3460
rect 4986 3414 5039 3426
rect -9283 2174 -9227 2186
rect -9283 2140 -9272 2174
rect -9238 2140 -9227 2174
rect -9283 2106 -9227 2140
rect -9283 2072 -9272 2106
rect -9238 2072 -9227 2106
rect -9283 2046 -9227 2072
rect -9107 2174 -9051 2186
rect -9107 2140 -9096 2174
rect -9062 2140 -9051 2174
rect -9107 2106 -9051 2140
rect -9107 2072 -9096 2106
rect -9062 2072 -9051 2106
rect -9107 2046 -9051 2072
rect -8931 2174 -8875 2186
rect -8931 2140 -8920 2174
rect -8886 2140 -8875 2174
rect -8931 2106 -8875 2140
rect -8931 2072 -8920 2106
rect -8886 2072 -8875 2106
rect -8931 2046 -8875 2072
rect -8755 2046 -8699 2186
rect -8579 2174 -8526 2186
rect -8579 2140 -8568 2174
rect -8534 2140 -8526 2174
rect -8579 2106 -8526 2140
rect -8579 2072 -8568 2106
rect -8534 2072 -8526 2106
rect -8579 2046 -8526 2072
<< mvpdiff >>
rect 3871 7152 3924 7170
rect 3871 7118 3879 7152
rect 3913 7118 3924 7152
rect 3871 7084 3924 7118
rect 3871 7050 3879 7084
rect 3913 7050 3924 7084
rect 3871 7016 3924 7050
rect 3871 6982 3879 7016
rect 3913 6982 3924 7016
rect 3871 6970 3924 6982
rect 4044 7152 4100 7170
rect 4044 7118 4055 7152
rect 4089 7118 4100 7152
rect 4044 7084 4100 7118
rect 4044 7050 4055 7084
rect 4089 7050 4100 7084
rect 4044 7016 4100 7050
rect 4044 6982 4055 7016
rect 4089 6982 4100 7016
rect 4044 6970 4100 6982
rect 4220 7152 4273 7170
rect 4220 7118 4231 7152
rect 4265 7118 4273 7152
rect 4220 7084 4273 7118
rect 4220 7050 4231 7084
rect 4265 7050 4273 7084
rect 4220 7016 4273 7050
rect 4220 6982 4231 7016
rect 4265 6982 4273 7016
rect 4220 6970 4273 6982
rect 4347 7152 4400 7170
rect 4347 7118 4355 7152
rect 4389 7118 4400 7152
rect 4347 7084 4400 7118
rect 4347 7050 4355 7084
rect 4389 7050 4400 7084
rect 4347 7016 4400 7050
rect 4347 6982 4355 7016
rect 4389 6982 4400 7016
rect 4347 6970 4400 6982
rect 4520 7152 4576 7170
rect 4520 7118 4531 7152
rect 4565 7118 4576 7152
rect 4520 7084 4576 7118
rect 4520 7050 4531 7084
rect 4565 7050 4576 7084
rect 4520 7016 4576 7050
rect 4520 6982 4531 7016
rect 4565 6982 4576 7016
rect 4520 6970 4576 6982
rect 4696 7152 4752 7170
rect 4696 7118 4707 7152
rect 4741 7118 4752 7152
rect 4696 7084 4752 7118
rect 4696 7050 4707 7084
rect 4741 7050 4752 7084
rect 4696 7016 4752 7050
rect 4696 6982 4707 7016
rect 4741 6982 4752 7016
rect 4696 6970 4752 6982
rect 4872 7152 4928 7170
rect 4872 7118 4883 7152
rect 4917 7118 4928 7152
rect 4872 7084 4928 7118
rect 4872 7050 4883 7084
rect 4917 7050 4928 7084
rect 4872 7016 4928 7050
rect 4872 6982 4883 7016
rect 4917 6982 4928 7016
rect 4872 6970 4928 6982
rect 5048 7152 5101 7170
rect 5048 7118 5059 7152
rect 5093 7118 5101 7152
rect 5048 7084 5101 7118
rect 5048 7050 5059 7084
rect 5093 7050 5101 7084
rect 5048 7016 5101 7050
rect 5048 6982 5059 7016
rect 5093 6982 5101 7016
rect 5048 6970 5101 6982
rect 5175 7152 5228 7170
rect 5175 7118 5183 7152
rect 5217 7118 5228 7152
rect 5175 7084 5228 7118
rect 5175 7050 5183 7084
rect 5217 7050 5228 7084
rect 5175 7016 5228 7050
rect 5175 6982 5183 7016
rect 5217 6982 5228 7016
rect 5175 6970 5228 6982
rect 5348 7152 5404 7170
rect 5348 7118 5359 7152
rect 5393 7118 5404 7152
rect 5348 7084 5404 7118
rect 5348 7050 5359 7084
rect 5393 7050 5404 7084
rect 5348 7016 5404 7050
rect 5348 6982 5359 7016
rect 5393 6982 5404 7016
rect 5348 6970 5404 6982
rect 5524 7152 5577 7170
rect 5524 7118 5535 7152
rect 5569 7118 5577 7152
rect 5524 7084 5577 7118
rect 5524 7050 5535 7084
rect 5569 7050 5577 7084
rect 5524 7016 5577 7050
rect 5524 6982 5535 7016
rect 5569 6982 5577 7016
rect 5524 6970 5577 6982
rect 5651 7152 5704 7170
rect 5651 7118 5659 7152
rect 5693 7118 5704 7152
rect 5651 7084 5704 7118
rect 5651 7050 5659 7084
rect 5693 7050 5704 7084
rect 5651 7016 5704 7050
rect 5651 6982 5659 7016
rect 5693 6982 5704 7016
rect 5651 6970 5704 6982
rect 5824 7152 5880 7170
rect 5824 7118 5835 7152
rect 5869 7118 5880 7152
rect 5824 7084 5880 7118
rect 5824 7050 5835 7084
rect 5869 7050 5880 7084
rect 5824 7016 5880 7050
rect 5824 6982 5835 7016
rect 5869 6982 5880 7016
rect 5824 6970 5880 6982
rect 6000 7152 6056 7170
rect 6000 7118 6011 7152
rect 6045 7118 6056 7152
rect 6000 7084 6056 7118
rect 6000 7050 6011 7084
rect 6045 7050 6056 7084
rect 6000 7016 6056 7050
rect 6000 6982 6011 7016
rect 6045 6982 6056 7016
rect 6000 6970 6056 6982
rect 6176 7152 6229 7170
rect 6176 7118 6187 7152
rect 6221 7118 6229 7152
rect 6176 7084 6229 7118
rect 6176 7050 6187 7084
rect 6221 7050 6229 7084
rect 6176 7016 6229 7050
rect 6176 6982 6187 7016
rect 6221 6982 6229 7016
rect 6176 6970 6229 6982
rect 3871 6890 3924 6902
rect 3871 6856 3879 6890
rect 3913 6856 3924 6890
rect 3871 6822 3924 6856
rect 3871 6788 3879 6822
rect 3913 6788 3924 6822
rect 3871 6754 3924 6788
rect 3871 6720 3879 6754
rect 3913 6720 3924 6754
rect 3871 6702 3924 6720
rect 4044 6890 4100 6902
rect 4044 6856 4055 6890
rect 4089 6856 4100 6890
rect 4044 6822 4100 6856
rect 4044 6788 4055 6822
rect 4089 6788 4100 6822
rect 4044 6754 4100 6788
rect 4044 6720 4055 6754
rect 4089 6720 4100 6754
rect 4044 6702 4100 6720
rect 4220 6890 4273 6902
rect 4220 6856 4231 6890
rect 4265 6856 4273 6890
rect 4220 6822 4273 6856
rect 4220 6788 4231 6822
rect 4265 6788 4273 6822
rect 4220 6754 4273 6788
rect 4220 6720 4231 6754
rect 4265 6720 4273 6754
rect 4220 6702 4273 6720
rect 4347 6890 4400 6902
rect 4347 6856 4355 6890
rect 4389 6856 4400 6890
rect 4347 6822 4400 6856
rect 4347 6788 4355 6822
rect 4389 6788 4400 6822
rect 4347 6754 4400 6788
rect 4347 6720 4355 6754
rect 4389 6720 4400 6754
rect 4347 6702 4400 6720
rect 4520 6890 4576 6902
rect 4520 6856 4531 6890
rect 4565 6856 4576 6890
rect 4520 6822 4576 6856
rect 4520 6788 4531 6822
rect 4565 6788 4576 6822
rect 4520 6754 4576 6788
rect 4520 6720 4531 6754
rect 4565 6720 4576 6754
rect 4520 6702 4576 6720
rect 4696 6890 4752 6902
rect 4696 6856 4707 6890
rect 4741 6856 4752 6890
rect 4696 6822 4752 6856
rect 4696 6788 4707 6822
rect 4741 6788 4752 6822
rect 4696 6754 4752 6788
rect 4696 6720 4707 6754
rect 4741 6720 4752 6754
rect 4696 6702 4752 6720
rect 4872 6890 4928 6902
rect 4872 6856 4883 6890
rect 4917 6856 4928 6890
rect 4872 6822 4928 6856
rect 4872 6788 4883 6822
rect 4917 6788 4928 6822
rect 4872 6754 4928 6788
rect 4872 6720 4883 6754
rect 4917 6720 4928 6754
rect 4872 6702 4928 6720
rect 5048 6890 5101 6902
rect 5048 6856 5059 6890
rect 5093 6856 5101 6890
rect 5048 6822 5101 6856
rect 5048 6788 5059 6822
rect 5093 6788 5101 6822
rect 5048 6754 5101 6788
rect 5048 6720 5059 6754
rect 5093 6720 5101 6754
rect 5048 6702 5101 6720
rect 5175 6890 5228 6902
rect 5175 6856 5183 6890
rect 5217 6856 5228 6890
rect 5175 6822 5228 6856
rect 5175 6788 5183 6822
rect 5217 6788 5228 6822
rect 5175 6754 5228 6788
rect 5175 6720 5183 6754
rect 5217 6720 5228 6754
rect 5175 6702 5228 6720
rect 5348 6890 5404 6902
rect 5348 6856 5359 6890
rect 5393 6856 5404 6890
rect 5348 6822 5404 6856
rect 5348 6788 5359 6822
rect 5393 6788 5404 6822
rect 5348 6754 5404 6788
rect 5348 6720 5359 6754
rect 5393 6720 5404 6754
rect 5348 6702 5404 6720
rect 5524 6890 5577 6902
rect 5524 6856 5535 6890
rect 5569 6856 5577 6890
rect 5524 6822 5577 6856
rect 5524 6788 5535 6822
rect 5569 6788 5577 6822
rect 5524 6754 5577 6788
rect 5524 6720 5535 6754
rect 5569 6720 5577 6754
rect 5524 6702 5577 6720
rect 5651 6890 5704 6902
rect 5651 6856 5659 6890
rect 5693 6856 5704 6890
rect 5651 6822 5704 6856
rect 5651 6788 5659 6822
rect 5693 6788 5704 6822
rect 5651 6754 5704 6788
rect 5651 6720 5659 6754
rect 5693 6720 5704 6754
rect 5651 6702 5704 6720
rect 5824 6890 5880 6902
rect 5824 6856 5835 6890
rect 5869 6856 5880 6890
rect 5824 6822 5880 6856
rect 5824 6788 5835 6822
rect 5869 6788 5880 6822
rect 5824 6754 5880 6788
rect 5824 6720 5835 6754
rect 5869 6720 5880 6754
rect 5824 6702 5880 6720
rect 6000 6890 6056 6902
rect 6000 6856 6011 6890
rect 6045 6856 6056 6890
rect 6000 6822 6056 6856
rect 6000 6788 6011 6822
rect 6045 6788 6056 6822
rect 6000 6754 6056 6788
rect 6000 6720 6011 6754
rect 6045 6720 6056 6754
rect 6000 6702 6056 6720
rect 6176 6890 6229 6902
rect 6176 6856 6187 6890
rect 6221 6856 6229 6890
rect 6176 6822 6229 6856
rect 6176 6788 6187 6822
rect 6221 6788 6229 6822
rect 6176 6754 6229 6788
rect 6176 6720 6187 6754
rect 6221 6720 6229 6754
rect 6176 6702 6229 6720
rect 3871 6516 3924 6534
rect 3871 6482 3879 6516
rect 3913 6482 3924 6516
rect 3871 6448 3924 6482
rect 3871 6414 3879 6448
rect 3913 6414 3924 6448
rect 3871 6380 3924 6414
rect 3871 6346 3879 6380
rect 3913 6346 3924 6380
rect 3871 6334 3924 6346
rect 4044 6516 4100 6534
rect 4044 6482 4055 6516
rect 4089 6482 4100 6516
rect 4044 6448 4100 6482
rect 4044 6414 4055 6448
rect 4089 6414 4100 6448
rect 4044 6380 4100 6414
rect 4044 6346 4055 6380
rect 4089 6346 4100 6380
rect 4044 6334 4100 6346
rect 4220 6516 4273 6534
rect 4220 6482 4231 6516
rect 4265 6482 4273 6516
rect 4220 6448 4273 6482
rect 4220 6414 4231 6448
rect 4265 6414 4273 6448
rect 4220 6380 4273 6414
rect 4220 6346 4231 6380
rect 4265 6346 4273 6380
rect 4220 6334 4273 6346
rect 4347 6516 4400 6534
rect 4347 6482 4355 6516
rect 4389 6482 4400 6516
rect 4347 6448 4400 6482
rect 4347 6414 4355 6448
rect 4389 6414 4400 6448
rect 4347 6380 4400 6414
rect 4347 6346 4355 6380
rect 4389 6346 4400 6380
rect 4347 6334 4400 6346
rect 4520 6516 4576 6534
rect 4520 6482 4531 6516
rect 4565 6482 4576 6516
rect 4520 6448 4576 6482
rect 4520 6414 4531 6448
rect 4565 6414 4576 6448
rect 4520 6380 4576 6414
rect 4520 6346 4531 6380
rect 4565 6346 4576 6380
rect 4520 6334 4576 6346
rect 4696 6516 4749 6534
rect 4696 6482 4707 6516
rect 4741 6482 4749 6516
rect 4696 6448 4749 6482
rect 4696 6414 4707 6448
rect 4741 6414 4749 6448
rect 4696 6380 4749 6414
rect 4696 6346 4707 6380
rect 4741 6346 4749 6380
rect 4696 6334 4749 6346
rect 4823 6516 4876 6534
rect 4823 6482 4831 6516
rect 4865 6482 4876 6516
rect 4823 6448 4876 6482
rect 4823 6414 4831 6448
rect 4865 6414 4876 6448
rect 4823 6380 4876 6414
rect 4823 6346 4831 6380
rect 4865 6346 4876 6380
rect 4823 6334 4876 6346
rect 4996 6516 5052 6534
rect 4996 6482 5007 6516
rect 5041 6482 5052 6516
rect 4996 6448 5052 6482
rect 4996 6414 5007 6448
rect 5041 6414 5052 6448
rect 4996 6380 5052 6414
rect 4996 6346 5007 6380
rect 5041 6346 5052 6380
rect 4996 6334 5052 6346
rect 5172 6516 5228 6534
rect 5172 6482 5183 6516
rect 5217 6482 5228 6516
rect 5172 6448 5228 6482
rect 5172 6414 5183 6448
rect 5217 6414 5228 6448
rect 5172 6380 5228 6414
rect 5172 6346 5183 6380
rect 5217 6346 5228 6380
rect 5172 6334 5228 6346
rect 5348 6516 5404 6534
rect 5348 6482 5359 6516
rect 5393 6482 5404 6516
rect 5348 6448 5404 6482
rect 5348 6414 5359 6448
rect 5393 6414 5404 6448
rect 5348 6380 5404 6414
rect 5348 6346 5359 6380
rect 5393 6346 5404 6380
rect 5348 6334 5404 6346
rect 5524 6516 5577 6534
rect 5524 6482 5535 6516
rect 5569 6482 5577 6516
rect 5524 6448 5577 6482
rect 5524 6414 5535 6448
rect 5569 6414 5577 6448
rect 5524 6380 5577 6414
rect 5524 6346 5535 6380
rect 5569 6346 5577 6380
rect 5524 6334 5577 6346
rect 5651 6516 5704 6534
rect 5651 6482 5659 6516
rect 5693 6482 5704 6516
rect 5651 6448 5704 6482
rect 5651 6414 5659 6448
rect 5693 6414 5704 6448
rect 5651 6380 5704 6414
rect 5651 6346 5659 6380
rect 5693 6346 5704 6380
rect 5651 6334 5704 6346
rect 5824 6516 5880 6534
rect 5824 6482 5835 6516
rect 5869 6482 5880 6516
rect 5824 6448 5880 6482
rect 5824 6414 5835 6448
rect 5869 6414 5880 6448
rect 5824 6380 5880 6414
rect 5824 6346 5835 6380
rect 5869 6346 5880 6380
rect 5824 6334 5880 6346
rect 6000 6516 6056 6534
rect 6000 6482 6011 6516
rect 6045 6482 6056 6516
rect 6000 6448 6056 6482
rect 6000 6414 6011 6448
rect 6045 6414 6056 6448
rect 6000 6380 6056 6414
rect 6000 6346 6011 6380
rect 6045 6346 6056 6380
rect 6000 6334 6056 6346
rect 6176 6516 6229 6534
rect 6176 6482 6187 6516
rect 6221 6482 6229 6516
rect 6176 6448 6229 6482
rect 6176 6414 6187 6448
rect 6221 6414 6229 6448
rect 6176 6380 6229 6414
rect 6176 6346 6187 6380
rect 6221 6346 6229 6380
rect 6176 6334 6229 6346
rect 3871 6254 3924 6266
rect 3871 6220 3879 6254
rect 3913 6220 3924 6254
rect 3871 6186 3924 6220
rect 3871 6152 3879 6186
rect 3913 6152 3924 6186
rect 3871 6118 3924 6152
rect 3871 6084 3879 6118
rect 3913 6084 3924 6118
rect 3871 6066 3924 6084
rect 4044 6254 4100 6266
rect 4044 6220 4055 6254
rect 4089 6220 4100 6254
rect 4044 6186 4100 6220
rect 4044 6152 4055 6186
rect 4089 6152 4100 6186
rect 4044 6066 4100 6152
rect 4220 6254 4273 6266
rect 4220 6220 4231 6254
rect 4265 6220 4273 6254
rect 4220 6186 4273 6220
rect 4220 6152 4231 6186
rect 4265 6152 4273 6186
rect 4220 6118 4273 6152
rect 4220 6084 4231 6118
rect 4265 6084 4273 6118
rect 4220 6066 4273 6084
rect 4347 6254 4400 6266
rect 4347 6220 4355 6254
rect 4389 6220 4400 6254
rect 4347 6186 4400 6220
rect 4347 6152 4355 6186
rect 4389 6152 4400 6186
rect 4347 6118 4400 6152
rect 4347 6084 4355 6118
rect 4389 6084 4400 6118
rect 4347 6066 4400 6084
rect 4520 6254 4576 6266
rect 4520 6220 4531 6254
rect 4565 6220 4576 6254
rect 4520 6186 4576 6220
rect 4520 6152 4531 6186
rect 4565 6152 4576 6186
rect 4520 6118 4576 6152
rect 4520 6084 4531 6118
rect 4565 6084 4576 6118
rect 4520 6066 4576 6084
rect 4696 6254 4749 6266
rect 4696 6220 4707 6254
rect 4741 6220 4749 6254
rect 4696 6186 4749 6220
rect 4696 6152 4707 6186
rect 4741 6152 4749 6186
rect 4696 6118 4749 6152
rect 4696 6084 4707 6118
rect 4741 6084 4749 6118
rect 4696 6066 4749 6084
rect 4823 6254 4876 6266
rect 4823 6220 4831 6254
rect 4865 6220 4876 6254
rect 4823 6186 4876 6220
rect 4823 6152 4831 6186
rect 4865 6152 4876 6186
rect 4823 6118 4876 6152
rect 4823 6084 4831 6118
rect 4865 6084 4876 6118
rect 4823 6066 4876 6084
rect 4996 6254 5052 6266
rect 4996 6220 5007 6254
rect 5041 6220 5052 6254
rect 4996 6186 5052 6220
rect 4996 6152 5007 6186
rect 5041 6152 5052 6186
rect 4996 6118 5052 6152
rect 4996 6084 5007 6118
rect 5041 6084 5052 6118
rect 4996 6066 5052 6084
rect 5172 6254 5228 6266
rect 5172 6220 5183 6254
rect 5217 6220 5228 6254
rect 5172 6186 5228 6220
rect 5172 6152 5183 6186
rect 5217 6152 5228 6186
rect 5172 6118 5228 6152
rect 5172 6084 5183 6118
rect 5217 6084 5228 6118
rect 5172 6066 5228 6084
rect 5348 6254 5404 6266
rect 5348 6220 5359 6254
rect 5393 6220 5404 6254
rect 5348 6186 5404 6220
rect 5348 6152 5359 6186
rect 5393 6152 5404 6186
rect 5348 6118 5404 6152
rect 5348 6084 5359 6118
rect 5393 6084 5404 6118
rect 5348 6066 5404 6084
rect 5524 6254 5577 6266
rect 5524 6220 5535 6254
rect 5569 6220 5577 6254
rect 5524 6186 5577 6220
rect 5524 6152 5535 6186
rect 5569 6152 5577 6186
rect 5524 6118 5577 6152
rect 5524 6084 5535 6118
rect 5569 6084 5577 6118
rect 5524 6066 5577 6084
rect 5651 6254 5704 6266
rect 5651 6220 5659 6254
rect 5693 6220 5704 6254
rect 5651 6186 5704 6220
rect 5651 6152 5659 6186
rect 5693 6152 5704 6186
rect 5651 6118 5704 6152
rect 5651 6084 5659 6118
rect 5693 6084 5704 6118
rect 5651 6066 5704 6084
rect 5824 6254 5880 6266
rect 5824 6220 5835 6254
rect 5869 6220 5880 6254
rect 5824 6186 5880 6220
rect 5824 6152 5835 6186
rect 5869 6152 5880 6186
rect 5824 6118 5880 6152
rect 5824 6084 5835 6118
rect 5869 6084 5880 6118
rect 5824 6066 5880 6084
rect 6000 6254 6056 6266
rect 6000 6220 6011 6254
rect 6045 6220 6056 6254
rect 6000 6186 6056 6220
rect 6000 6152 6011 6186
rect 6045 6152 6056 6186
rect 6000 6118 6056 6152
rect 6000 6084 6011 6118
rect 6045 6084 6056 6118
rect 6000 6066 6056 6084
rect 6176 6254 6229 6266
rect 6176 6220 6187 6254
rect 6221 6220 6229 6254
rect 6176 6186 6229 6220
rect 6176 6152 6187 6186
rect 6221 6152 6229 6186
rect 6176 6118 6229 6152
rect 6176 6084 6187 6118
rect 6221 6084 6229 6118
rect 6176 6066 6229 6084
rect 3966 5075 4019 5087
rect 3966 5041 3974 5075
rect 4008 5041 4019 5075
rect 3966 5007 4019 5041
rect 3966 4973 3974 5007
rect 4008 4973 4019 5007
rect 3966 4939 4019 4973
rect 3966 4905 3974 4939
rect 4008 4905 4019 4939
rect 3966 4887 4019 4905
rect 4139 5075 4195 5087
rect 4139 5041 4150 5075
rect 4184 5041 4195 5075
rect 4139 5007 4195 5041
rect 4139 4973 4150 5007
rect 4184 4973 4195 5007
rect 4139 4939 4195 4973
rect 4139 4905 4150 4939
rect 4184 4905 4195 4939
rect 4139 4887 4195 4905
rect 4315 5075 4371 5087
rect 4315 5041 4326 5075
rect 4360 5041 4371 5075
rect 4315 5007 4371 5041
rect 4315 4973 4326 5007
rect 4360 4973 4371 5007
rect 4315 4939 4371 4973
rect 4315 4905 4326 4939
rect 4360 4905 4371 4939
rect 4315 4887 4371 4905
rect 4491 5075 4547 5087
rect 4491 5041 4502 5075
rect 4536 5041 4547 5075
rect 4491 5007 4547 5041
rect 4491 4973 4502 5007
rect 4536 4973 4547 5007
rect 4491 4939 4547 4973
rect 4491 4905 4502 4939
rect 4536 4905 4547 4939
rect 4491 4887 4547 4905
rect 4667 5075 4723 5087
rect 4667 5041 4678 5075
rect 4712 5041 4723 5075
rect 4667 5007 4723 5041
rect 4667 4973 4678 5007
rect 4712 4973 4723 5007
rect 4667 4939 4723 4973
rect 4667 4905 4678 4939
rect 4712 4905 4723 4939
rect 4667 4887 4723 4905
rect 4843 5075 4899 5087
rect 4843 5041 4854 5075
rect 4888 5041 4899 5075
rect 4843 5007 4899 5041
rect 4843 4973 4854 5007
rect 4888 4973 4899 5007
rect 4843 4939 4899 4973
rect 4843 4905 4854 4939
rect 4888 4905 4899 4939
rect 4843 4887 4899 4905
rect 5019 5075 5072 5087
rect 5019 5041 5030 5075
rect 5064 5041 5072 5075
rect 5019 5007 5072 5041
rect 5019 4973 5030 5007
rect 5064 4973 5072 5007
rect 5019 4939 5072 4973
rect 5019 4905 5030 4939
rect 5064 4905 5072 4939
rect 5019 4887 5072 4905
rect 5340 5026 5393 5044
rect 5340 4992 5348 5026
rect 5382 4992 5393 5026
rect 5340 4958 5393 4992
rect 5340 4924 5348 4958
rect 5382 4924 5393 4958
rect 5340 4890 5393 4924
rect 5340 4856 5348 4890
rect 5382 4856 5393 4890
rect 5340 4844 5393 4856
rect 5513 5026 5566 5044
rect 5513 4992 5524 5026
rect 5558 4992 5566 5026
rect 5513 4958 5566 4992
rect 5513 4924 5524 4958
rect 5558 4924 5566 4958
rect 5513 4890 5566 4924
rect 5513 4856 5524 4890
rect 5558 4856 5566 4890
rect 5513 4844 5566 4856
rect 5640 5026 5693 5044
rect 5640 4992 5648 5026
rect 5682 4992 5693 5026
rect 5640 4958 5693 4992
rect 5640 4924 5648 4958
rect 5682 4924 5693 4958
rect 5640 4890 5693 4924
rect 5640 4856 5648 4890
rect 5682 4856 5693 4890
rect 5640 4844 5693 4856
rect 5813 5026 5869 5044
rect 5813 4992 5824 5026
rect 5858 4992 5869 5026
rect 5813 4958 5869 4992
rect 5813 4924 5824 4958
rect 5858 4924 5869 4958
rect 5813 4890 5869 4924
rect 5813 4856 5824 4890
rect 5858 4856 5869 4890
rect 5813 4844 5869 4856
rect 5989 5026 6045 5044
rect 5989 4992 6000 5026
rect 6034 4992 6045 5026
rect 5989 4958 6045 4992
rect 5989 4924 6000 4958
rect 6034 4924 6045 4958
rect 5989 4890 6045 4924
rect 5989 4856 6000 4890
rect 6034 4856 6045 4890
rect 5989 4844 6045 4856
rect 6165 5026 6218 5044
rect 6165 4992 6176 5026
rect 6210 4992 6218 5026
rect 6165 4958 6218 4992
rect 6165 4924 6176 4958
rect 6210 4924 6218 4958
rect 6165 4890 6218 4924
rect 6165 4856 6176 4890
rect 6210 4856 6218 4890
rect 6165 4844 6218 4856
rect 3966 4807 4019 4819
rect 3966 4773 3974 4807
rect 4008 4773 4019 4807
rect 3966 4739 4019 4773
rect 3966 4705 3974 4739
rect 4008 4705 4019 4739
rect 3966 4671 4019 4705
rect 3966 4637 3974 4671
rect 4008 4637 4019 4671
rect 3966 4619 4019 4637
rect 4139 4807 4195 4819
rect 4139 4773 4150 4807
rect 4184 4773 4195 4807
rect 4139 4739 4195 4773
rect 4139 4705 4150 4739
rect 4184 4705 4195 4739
rect 4139 4671 4195 4705
rect 4139 4637 4150 4671
rect 4184 4637 4195 4671
rect 4139 4619 4195 4637
rect 4315 4807 4371 4819
rect 4315 4773 4326 4807
rect 4360 4773 4371 4807
rect 4315 4739 4371 4773
rect 4315 4705 4326 4739
rect 4360 4705 4371 4739
rect 4315 4671 4371 4705
rect 4315 4637 4326 4671
rect 4360 4637 4371 4671
rect 4315 4619 4371 4637
rect 4491 4807 4547 4819
rect 4491 4773 4502 4807
rect 4536 4773 4547 4807
rect 4491 4739 4547 4773
rect 4491 4705 4502 4739
rect 4536 4705 4547 4739
rect 4491 4671 4547 4705
rect 4491 4637 4502 4671
rect 4536 4637 4547 4671
rect 4491 4619 4547 4637
rect 4667 4807 4723 4819
rect 4667 4773 4678 4807
rect 4712 4773 4723 4807
rect 4667 4739 4723 4773
rect 4667 4705 4678 4739
rect 4712 4705 4723 4739
rect 4667 4671 4723 4705
rect 4667 4637 4678 4671
rect 4712 4637 4723 4671
rect 4667 4619 4723 4637
rect 4843 4807 4899 4819
rect 4843 4773 4854 4807
rect 4888 4773 4899 4807
rect 4843 4739 4899 4773
rect 4843 4705 4854 4739
rect 4888 4705 4899 4739
rect 4843 4671 4899 4705
rect 4843 4637 4854 4671
rect 4888 4637 4899 4671
rect 4843 4619 4899 4637
rect 5019 4807 5072 4819
rect 5019 4773 5030 4807
rect 5064 4773 5072 4807
rect 5019 4739 5072 4773
rect 5019 4705 5030 4739
rect 5064 4705 5072 4739
rect 5019 4671 5072 4705
rect 5019 4637 5030 4671
rect 5064 4637 5072 4671
rect 5019 4619 5072 4637
rect 5340 4764 5393 4776
rect 5340 4730 5348 4764
rect 5382 4730 5393 4764
rect 5340 4696 5393 4730
rect 5340 4662 5348 4696
rect 5382 4662 5393 4696
rect 5340 4628 5393 4662
rect 5340 4594 5348 4628
rect 5382 4594 5393 4628
rect 5340 4576 5393 4594
rect 5513 4764 5566 4776
rect 5513 4730 5524 4764
rect 5558 4730 5566 4764
rect 5513 4696 5566 4730
rect 5513 4662 5524 4696
rect 5558 4662 5566 4696
rect 5513 4628 5566 4662
rect 5513 4594 5524 4628
rect 5558 4594 5566 4628
rect 5513 4576 5566 4594
rect 5640 4764 5693 4776
rect 5640 4730 5648 4764
rect 5682 4730 5693 4764
rect 5640 4696 5693 4730
rect 5640 4662 5648 4696
rect 5682 4662 5693 4696
rect 5640 4628 5693 4662
rect 5640 4594 5648 4628
rect 5682 4594 5693 4628
rect 5640 4576 5693 4594
rect 5813 4764 5869 4776
rect 5813 4730 5824 4764
rect 5858 4730 5869 4764
rect 5813 4696 5869 4730
rect 5813 4662 5824 4696
rect 5858 4662 5869 4696
rect 5813 4628 5869 4662
rect 5813 4594 5824 4628
rect 5858 4594 5869 4628
rect 5813 4576 5869 4594
rect 5989 4764 6045 4776
rect 5989 4730 6000 4764
rect 6034 4730 6045 4764
rect 5989 4696 6045 4730
rect 5989 4662 6000 4696
rect 6034 4662 6045 4696
rect 5989 4628 6045 4662
rect 5989 4594 6000 4628
rect 6034 4594 6045 4628
rect 5989 4576 6045 4594
rect 6165 4764 6218 4776
rect 6165 4730 6176 4764
rect 6210 4730 6218 4764
rect 6165 4696 6218 4730
rect 6165 4662 6176 4696
rect 6210 4662 6218 4696
rect 6165 4628 6218 4662
rect 6165 4594 6176 4628
rect 6210 4594 6218 4628
rect 6165 4576 6218 4594
rect 5315 4374 5368 4392
rect 5315 4340 5323 4374
rect 5357 4340 5368 4374
rect 5315 4306 5368 4340
rect 3933 4266 3986 4284
rect 3933 4232 3941 4266
rect 3975 4232 3986 4266
rect 3933 4198 3986 4232
rect 3933 4164 3941 4198
rect 3975 4164 3986 4198
rect 3933 4130 3986 4164
rect 3933 4096 3941 4130
rect 3975 4096 3986 4130
rect 3933 4084 3986 4096
rect 4106 4266 4162 4284
rect 4106 4232 4117 4266
rect 4151 4232 4162 4266
rect 4106 4198 4162 4232
rect 4106 4164 4117 4198
rect 4151 4164 4162 4198
rect 4106 4130 4162 4164
rect 4106 4096 4117 4130
rect 4151 4096 4162 4130
rect 4106 4084 4162 4096
rect 4282 4266 4338 4284
rect 4282 4232 4293 4266
rect 4327 4232 4338 4266
rect 4282 4198 4338 4232
rect 4282 4164 4293 4198
rect 4327 4164 4338 4198
rect 4282 4130 4338 4164
rect 4282 4096 4293 4130
rect 4327 4096 4338 4130
rect 4282 4084 4338 4096
rect 4458 4266 4514 4284
rect 4458 4232 4469 4266
rect 4503 4232 4514 4266
rect 4458 4198 4514 4232
rect 4458 4164 4469 4198
rect 4503 4164 4514 4198
rect 4458 4130 4514 4164
rect 4458 4096 4469 4130
rect 4503 4096 4514 4130
rect 4458 4084 4514 4096
rect 4634 4266 4690 4284
rect 4634 4232 4645 4266
rect 4679 4232 4690 4266
rect 4634 4198 4690 4232
rect 4634 4164 4645 4198
rect 4679 4164 4690 4198
rect 4634 4130 4690 4164
rect 4634 4096 4645 4130
rect 4679 4096 4690 4130
rect 4634 4084 4690 4096
rect 4810 4266 4866 4284
rect 4810 4232 4821 4266
rect 4855 4232 4866 4266
rect 4810 4198 4866 4232
rect 4810 4164 4821 4198
rect 4855 4164 4866 4198
rect 4810 4130 4866 4164
rect 4810 4096 4821 4130
rect 4855 4096 4866 4130
rect 4810 4084 4866 4096
rect 4986 4266 5039 4284
rect 4986 4232 4997 4266
rect 5031 4232 5039 4266
rect 4986 4198 5039 4232
rect 4986 4164 4997 4198
rect 5031 4164 5039 4198
rect 5315 4272 5323 4306
rect 5357 4272 5368 4306
rect 5315 4238 5368 4272
rect 5315 4204 5323 4238
rect 5357 4204 5368 4238
rect 5315 4192 5368 4204
rect 5488 4374 5544 4392
rect 5488 4340 5499 4374
rect 5533 4340 5544 4374
rect 5488 4306 5544 4340
rect 5488 4272 5499 4306
rect 5533 4272 5544 4306
rect 5488 4238 5544 4272
rect 5488 4204 5499 4238
rect 5533 4204 5544 4238
rect 5488 4192 5544 4204
rect 5664 4374 5720 4392
rect 5664 4340 5675 4374
rect 5709 4340 5720 4374
rect 5664 4306 5720 4340
rect 5664 4272 5675 4306
rect 5709 4272 5720 4306
rect 5664 4238 5720 4272
rect 5664 4204 5675 4238
rect 5709 4204 5720 4238
rect 5664 4192 5720 4204
rect 5840 4374 5896 4392
rect 5840 4340 5851 4374
rect 5885 4340 5896 4374
rect 5840 4306 5896 4340
rect 5840 4272 5851 4306
rect 5885 4272 5896 4306
rect 5840 4238 5896 4272
rect 5840 4204 5851 4238
rect 5885 4204 5896 4238
rect 5840 4192 5896 4204
rect 6016 4374 6072 4392
rect 6016 4340 6027 4374
rect 6061 4340 6072 4374
rect 6016 4306 6072 4340
rect 6016 4272 6027 4306
rect 6061 4272 6072 4306
rect 6016 4238 6072 4272
rect 6016 4204 6027 4238
rect 6061 4204 6072 4238
rect 6016 4192 6072 4204
rect 6192 4374 6245 4392
rect 6192 4340 6203 4374
rect 6237 4340 6245 4374
rect 6192 4306 6245 4340
rect 6192 4272 6203 4306
rect 6237 4272 6245 4306
rect 6192 4238 6245 4272
rect 6192 4204 6203 4238
rect 6237 4204 6245 4238
rect 6192 4192 6245 4204
rect 4986 4130 5039 4164
rect 4986 4096 4997 4130
rect 5031 4096 5039 4130
rect 4986 4084 5039 4096
rect 5315 4112 5368 4124
rect 5315 4078 5323 4112
rect 5357 4078 5368 4112
rect 5315 4044 5368 4078
rect 3933 3998 3986 4016
rect 3933 3964 3941 3998
rect 3975 3964 3986 3998
rect 3933 3930 3986 3964
rect 3933 3896 3941 3930
rect 3975 3896 3986 3930
rect 3933 3862 3986 3896
rect 3933 3828 3941 3862
rect 3975 3828 3986 3862
rect 3933 3816 3986 3828
rect 4106 3998 4162 4016
rect 4106 3964 4117 3998
rect 4151 3964 4162 3998
rect 4106 3930 4162 3964
rect 4106 3896 4117 3930
rect 4151 3896 4162 3930
rect 4106 3862 4162 3896
rect 4106 3828 4117 3862
rect 4151 3828 4162 3862
rect 4106 3816 4162 3828
rect 4282 3998 4338 4016
rect 4282 3964 4293 3998
rect 4327 3964 4338 3998
rect 4282 3930 4338 3964
rect 4282 3896 4293 3930
rect 4327 3896 4338 3930
rect 4282 3862 4338 3896
rect 4282 3828 4293 3862
rect 4327 3828 4338 3862
rect 4282 3816 4338 3828
rect 4458 3998 4514 4016
rect 4458 3964 4469 3998
rect 4503 3964 4514 3998
rect 4458 3930 4514 3964
rect 4458 3896 4469 3930
rect 4503 3896 4514 3930
rect 4458 3862 4514 3896
rect 4458 3828 4469 3862
rect 4503 3828 4514 3862
rect 4458 3816 4514 3828
rect 4634 3998 4690 4016
rect 4634 3964 4645 3998
rect 4679 3964 4690 3998
rect 4634 3930 4690 3964
rect 4634 3896 4645 3930
rect 4679 3896 4690 3930
rect 4634 3862 4690 3896
rect 4634 3828 4645 3862
rect 4679 3828 4690 3862
rect 4634 3816 4690 3828
rect 4810 3998 4866 4016
rect 4810 3964 4821 3998
rect 4855 3964 4866 3998
rect 4810 3930 4866 3964
rect 4810 3896 4821 3930
rect 4855 3896 4866 3930
rect 4810 3862 4866 3896
rect 4810 3828 4821 3862
rect 4855 3828 4866 3862
rect 4810 3816 4866 3828
rect 4986 3998 5039 4016
rect 4986 3964 4997 3998
rect 5031 3964 5039 3998
rect 4986 3930 5039 3964
rect 4986 3896 4997 3930
rect 5031 3896 5039 3930
rect 5315 4010 5323 4044
rect 5357 4010 5368 4044
rect 5315 3976 5368 4010
rect 5315 3942 5323 3976
rect 5357 3942 5368 3976
rect 5315 3924 5368 3942
rect 5488 4112 5544 4124
rect 5488 4078 5499 4112
rect 5533 4078 5544 4112
rect 5488 4044 5544 4078
rect 5488 4010 5499 4044
rect 5533 4010 5544 4044
rect 5488 3924 5544 4010
rect 5664 4112 5720 4124
rect 5664 4078 5675 4112
rect 5709 4078 5720 4112
rect 5664 4044 5720 4078
rect 5664 4010 5675 4044
rect 5709 4010 5720 4044
rect 5664 3976 5720 4010
rect 5664 3942 5675 3976
rect 5709 3942 5720 3976
rect 5664 3924 5720 3942
rect 5840 4112 5896 4124
rect 5840 4078 5851 4112
rect 5885 4078 5896 4112
rect 5840 4044 5896 4078
rect 5840 4010 5851 4044
rect 5885 4010 5896 4044
rect 5840 3976 5896 4010
rect 5840 3942 5851 3976
rect 5885 3942 5896 3976
rect 5840 3924 5896 3942
rect 6016 4112 6072 4124
rect 6016 4078 6027 4112
rect 6061 4078 6072 4112
rect 6016 4044 6072 4078
rect 6016 4010 6027 4044
rect 6061 4010 6072 4044
rect 6016 3976 6072 4010
rect 6016 3942 6027 3976
rect 6061 3942 6072 3976
rect 6016 3924 6072 3942
rect 6192 4112 6245 4124
rect 6192 4078 6203 4112
rect 6237 4078 6245 4112
rect 6192 4044 6245 4078
rect 6192 4010 6203 4044
rect 6237 4010 6245 4044
rect 6192 3976 6245 4010
rect 6192 3942 6203 3976
rect 6237 3942 6245 3976
rect 6192 3924 6245 3942
rect 4986 3862 5039 3896
rect 4986 3828 4997 3862
rect 5031 3828 5039 3862
rect 4986 3816 5039 3828
rect -9280 2834 -9227 2852
rect -9280 2800 -9272 2834
rect -9238 2800 -9227 2834
rect -9280 2766 -9227 2800
rect -9280 2732 -9272 2766
rect -9238 2732 -9227 2766
rect -9280 2698 -9227 2732
rect -9280 2664 -9272 2698
rect -9238 2664 -9227 2698
rect -9280 2652 -9227 2664
rect -9107 2834 -9051 2852
rect -9107 2800 -9096 2834
rect -9062 2800 -9051 2834
rect -9107 2766 -9051 2800
rect -9107 2732 -9096 2766
rect -9062 2732 -9051 2766
rect -9107 2698 -9051 2732
rect -9107 2664 -9096 2698
rect -9062 2664 -9051 2698
rect -9107 2652 -9051 2664
rect -8931 2834 -8875 2852
rect -8931 2800 -8920 2834
rect -8886 2800 -8875 2834
rect -8931 2766 -8875 2800
rect -8931 2732 -8920 2766
rect -8886 2732 -8875 2766
rect -8931 2698 -8875 2732
rect -8931 2664 -8920 2698
rect -8886 2664 -8875 2698
rect -8931 2652 -8875 2664
rect -8755 2834 -8699 2852
rect -8755 2800 -8744 2834
rect -8710 2800 -8699 2834
rect -8755 2766 -8699 2800
rect -8755 2732 -8744 2766
rect -8710 2732 -8699 2766
rect -8755 2698 -8699 2732
rect -8755 2664 -8744 2698
rect -8710 2664 -8699 2698
rect -8755 2652 -8699 2664
rect -8579 2834 -8526 2852
rect -8579 2800 -8568 2834
rect -8534 2800 -8526 2834
rect -8579 2766 -8526 2800
rect -8579 2732 -8568 2766
rect -8534 2732 -8526 2766
rect -8579 2698 -8526 2732
rect -8579 2664 -8568 2698
rect -8534 2664 -8526 2698
rect -8579 2652 -8526 2664
rect -9280 2572 -9227 2584
rect -9280 2538 -9272 2572
rect -9238 2538 -9227 2572
rect -9280 2504 -9227 2538
rect -9280 2470 -9272 2504
rect -9238 2470 -9227 2504
rect -9280 2436 -9227 2470
rect -9280 2402 -9272 2436
rect -9238 2402 -9227 2436
rect -9280 2384 -9227 2402
rect -9107 2572 -9051 2584
rect -9107 2538 -9096 2572
rect -9062 2538 -9051 2572
rect -9107 2504 -9051 2538
rect -9107 2470 -9096 2504
rect -9062 2470 -9051 2504
rect -9107 2384 -9051 2470
rect -8931 2572 -8875 2584
rect -8931 2538 -8920 2572
rect -8886 2538 -8875 2572
rect -8931 2504 -8875 2538
rect -8931 2470 -8920 2504
rect -8886 2470 -8875 2504
rect -8931 2436 -8875 2470
rect -8931 2402 -8920 2436
rect -8886 2402 -8875 2436
rect -8931 2384 -8875 2402
rect -8755 2572 -8699 2584
rect -8755 2538 -8744 2572
rect -8710 2538 -8699 2572
rect -8755 2504 -8699 2538
rect -8755 2470 -8744 2504
rect -8710 2470 -8699 2504
rect -8755 2436 -8699 2470
rect -8755 2402 -8744 2436
rect -8710 2402 -8699 2436
rect -8755 2384 -8699 2402
rect -8579 2572 -8526 2584
rect -8579 2538 -8568 2572
rect -8534 2538 -8526 2572
rect -8579 2504 -8526 2538
rect -8579 2470 -8568 2504
rect -8534 2470 -8526 2504
rect -8579 2436 -8526 2470
rect -8579 2402 -8568 2436
rect -8534 2402 -8526 2436
rect -8579 2384 -8526 2402
<< mvndiffc >>
rect 3879 7448 3913 7482
rect 3879 7380 3913 7414
rect 4231 7448 4265 7482
rect 4231 7380 4265 7414
rect 4355 7448 4389 7482
rect 4355 7380 4389 7414
rect 4707 7448 4741 7482
rect 4707 7380 4741 7414
rect 5059 7448 5093 7482
rect 5059 7380 5093 7414
rect 5183 7448 5217 7482
rect 5183 7380 5217 7414
rect 5535 7448 5569 7482
rect 5535 7380 5569 7414
rect 5659 7448 5693 7482
rect 5659 7380 5693 7414
rect 5835 7448 5869 7482
rect 5835 7380 5869 7414
rect 6011 7448 6045 7482
rect 6011 7380 6045 7414
rect 6187 7448 6221 7482
rect 6187 7380 6221 7414
rect 3879 5822 3913 5856
rect 3879 5754 3913 5788
rect 4055 5822 4089 5856
rect 4055 5754 4089 5788
rect 4231 5822 4265 5856
rect 4231 5754 4265 5788
rect 4355 5822 4389 5856
rect 4355 5754 4389 5788
rect 4707 5822 4741 5856
rect 4707 5754 4741 5788
rect 4831 5822 4865 5856
rect 4831 5754 4865 5788
rect 5183 5822 5217 5856
rect 5183 5754 5217 5788
rect 5535 5822 5569 5856
rect 5535 5754 5569 5788
rect 5659 5822 5693 5856
rect 5659 5754 5693 5788
rect 5835 5822 5869 5856
rect 5835 5754 5869 5788
rect 6011 5822 6045 5856
rect 6011 5754 6045 5788
rect 6187 5822 6221 5856
rect 6187 5754 6221 5788
rect 3974 5443 4008 5477
rect 3974 5375 4008 5409
rect 4150 5443 4184 5477
rect 4150 5375 4184 5409
rect 4326 5443 4360 5477
rect 4326 5375 4360 5409
rect 4502 5443 4536 5477
rect 4502 5375 4536 5409
rect 4678 5443 4712 5477
rect 4678 5375 4712 5409
rect 4854 5443 4888 5477
rect 4854 5375 4888 5409
rect 5030 5443 5064 5477
rect 5030 5375 5064 5409
rect 5348 5322 5382 5356
rect 5348 5254 5382 5288
rect 5524 5322 5558 5356
rect 5524 5254 5558 5288
rect 5648 5322 5682 5356
rect 5648 5254 5682 5288
rect 5824 5322 5858 5356
rect 5824 5254 5858 5288
rect 6000 5322 6034 5356
rect 6000 5254 6034 5288
rect 6176 5322 6210 5356
rect 6176 5254 6210 5288
rect 5323 3680 5357 3714
rect 5323 3612 5357 3646
rect 5499 3680 5533 3714
rect 5499 3612 5533 3646
rect 5675 3680 5709 3714
rect 5675 3612 5709 3646
rect 5851 3680 5885 3714
rect 5851 3612 5885 3646
rect 6027 3680 6061 3714
rect 6027 3612 6061 3646
rect 6203 3680 6237 3714
rect 6203 3612 6237 3646
rect 3941 3494 3975 3528
rect 3941 3426 3975 3460
rect 4117 3494 4151 3528
rect 4117 3426 4151 3460
rect 4293 3494 4327 3528
rect 4293 3426 4327 3460
rect 4469 3494 4503 3528
rect 4469 3426 4503 3460
rect 4645 3494 4679 3528
rect 4645 3426 4679 3460
rect 4821 3494 4855 3528
rect 4821 3426 4855 3460
rect 4997 3494 5031 3528
rect 4997 3426 5031 3460
rect -9272 2140 -9238 2174
rect -9272 2072 -9238 2106
rect -9096 2140 -9062 2174
rect -9096 2072 -9062 2106
rect -8920 2140 -8886 2174
rect -8920 2072 -8886 2106
rect -8568 2140 -8534 2174
rect -8568 2072 -8534 2106
<< mvpdiffc >>
rect 3879 7118 3913 7152
rect 3879 7050 3913 7084
rect 3879 6982 3913 7016
rect 4055 7118 4089 7152
rect 4055 7050 4089 7084
rect 4055 6982 4089 7016
rect 4231 7118 4265 7152
rect 4231 7050 4265 7084
rect 4231 6982 4265 7016
rect 4355 7118 4389 7152
rect 4355 7050 4389 7084
rect 4355 6982 4389 7016
rect 4531 7118 4565 7152
rect 4531 7050 4565 7084
rect 4531 6982 4565 7016
rect 4707 7118 4741 7152
rect 4707 7050 4741 7084
rect 4707 6982 4741 7016
rect 4883 7118 4917 7152
rect 4883 7050 4917 7084
rect 4883 6982 4917 7016
rect 5059 7118 5093 7152
rect 5059 7050 5093 7084
rect 5059 6982 5093 7016
rect 5183 7118 5217 7152
rect 5183 7050 5217 7084
rect 5183 6982 5217 7016
rect 5359 7118 5393 7152
rect 5359 7050 5393 7084
rect 5359 6982 5393 7016
rect 5535 7118 5569 7152
rect 5535 7050 5569 7084
rect 5535 6982 5569 7016
rect 5659 7118 5693 7152
rect 5659 7050 5693 7084
rect 5659 6982 5693 7016
rect 5835 7118 5869 7152
rect 5835 7050 5869 7084
rect 5835 6982 5869 7016
rect 6011 7118 6045 7152
rect 6011 7050 6045 7084
rect 6011 6982 6045 7016
rect 6187 7118 6221 7152
rect 6187 7050 6221 7084
rect 6187 6982 6221 7016
rect 3879 6856 3913 6890
rect 3879 6788 3913 6822
rect 3879 6720 3913 6754
rect 4055 6856 4089 6890
rect 4055 6788 4089 6822
rect 4055 6720 4089 6754
rect 4231 6856 4265 6890
rect 4231 6788 4265 6822
rect 4231 6720 4265 6754
rect 4355 6856 4389 6890
rect 4355 6788 4389 6822
rect 4355 6720 4389 6754
rect 4531 6856 4565 6890
rect 4531 6788 4565 6822
rect 4531 6720 4565 6754
rect 4707 6856 4741 6890
rect 4707 6788 4741 6822
rect 4707 6720 4741 6754
rect 4883 6856 4917 6890
rect 4883 6788 4917 6822
rect 4883 6720 4917 6754
rect 5059 6856 5093 6890
rect 5059 6788 5093 6822
rect 5059 6720 5093 6754
rect 5183 6856 5217 6890
rect 5183 6788 5217 6822
rect 5183 6720 5217 6754
rect 5359 6856 5393 6890
rect 5359 6788 5393 6822
rect 5359 6720 5393 6754
rect 5535 6856 5569 6890
rect 5535 6788 5569 6822
rect 5535 6720 5569 6754
rect 5659 6856 5693 6890
rect 5659 6788 5693 6822
rect 5659 6720 5693 6754
rect 5835 6856 5869 6890
rect 5835 6788 5869 6822
rect 5835 6720 5869 6754
rect 6011 6856 6045 6890
rect 6011 6788 6045 6822
rect 6011 6720 6045 6754
rect 6187 6856 6221 6890
rect 6187 6788 6221 6822
rect 6187 6720 6221 6754
rect 3879 6482 3913 6516
rect 3879 6414 3913 6448
rect 3879 6346 3913 6380
rect 4055 6482 4089 6516
rect 4055 6414 4089 6448
rect 4055 6346 4089 6380
rect 4231 6482 4265 6516
rect 4231 6414 4265 6448
rect 4231 6346 4265 6380
rect 4355 6482 4389 6516
rect 4355 6414 4389 6448
rect 4355 6346 4389 6380
rect 4531 6482 4565 6516
rect 4531 6414 4565 6448
rect 4531 6346 4565 6380
rect 4707 6482 4741 6516
rect 4707 6414 4741 6448
rect 4707 6346 4741 6380
rect 4831 6482 4865 6516
rect 4831 6414 4865 6448
rect 4831 6346 4865 6380
rect 5007 6482 5041 6516
rect 5007 6414 5041 6448
rect 5007 6346 5041 6380
rect 5183 6482 5217 6516
rect 5183 6414 5217 6448
rect 5183 6346 5217 6380
rect 5359 6482 5393 6516
rect 5359 6414 5393 6448
rect 5359 6346 5393 6380
rect 5535 6482 5569 6516
rect 5535 6414 5569 6448
rect 5535 6346 5569 6380
rect 5659 6482 5693 6516
rect 5659 6414 5693 6448
rect 5659 6346 5693 6380
rect 5835 6482 5869 6516
rect 5835 6414 5869 6448
rect 5835 6346 5869 6380
rect 6011 6482 6045 6516
rect 6011 6414 6045 6448
rect 6011 6346 6045 6380
rect 6187 6482 6221 6516
rect 6187 6414 6221 6448
rect 6187 6346 6221 6380
rect 3879 6220 3913 6254
rect 3879 6152 3913 6186
rect 3879 6084 3913 6118
rect 4055 6220 4089 6254
rect 4055 6152 4089 6186
rect 4231 6220 4265 6254
rect 4231 6152 4265 6186
rect 4231 6084 4265 6118
rect 4355 6220 4389 6254
rect 4355 6152 4389 6186
rect 4355 6084 4389 6118
rect 4531 6220 4565 6254
rect 4531 6152 4565 6186
rect 4531 6084 4565 6118
rect 4707 6220 4741 6254
rect 4707 6152 4741 6186
rect 4707 6084 4741 6118
rect 4831 6220 4865 6254
rect 4831 6152 4865 6186
rect 4831 6084 4865 6118
rect 5007 6220 5041 6254
rect 5007 6152 5041 6186
rect 5007 6084 5041 6118
rect 5183 6220 5217 6254
rect 5183 6152 5217 6186
rect 5183 6084 5217 6118
rect 5359 6220 5393 6254
rect 5359 6152 5393 6186
rect 5359 6084 5393 6118
rect 5535 6220 5569 6254
rect 5535 6152 5569 6186
rect 5535 6084 5569 6118
rect 5659 6220 5693 6254
rect 5659 6152 5693 6186
rect 5659 6084 5693 6118
rect 5835 6220 5869 6254
rect 5835 6152 5869 6186
rect 5835 6084 5869 6118
rect 6011 6220 6045 6254
rect 6011 6152 6045 6186
rect 6011 6084 6045 6118
rect 6187 6220 6221 6254
rect 6187 6152 6221 6186
rect 6187 6084 6221 6118
rect 3974 5041 4008 5075
rect 3974 4973 4008 5007
rect 3974 4905 4008 4939
rect 4150 5041 4184 5075
rect 4150 4973 4184 5007
rect 4150 4905 4184 4939
rect 4326 5041 4360 5075
rect 4326 4973 4360 5007
rect 4326 4905 4360 4939
rect 4502 5041 4536 5075
rect 4502 4973 4536 5007
rect 4502 4905 4536 4939
rect 4678 5041 4712 5075
rect 4678 4973 4712 5007
rect 4678 4905 4712 4939
rect 4854 5041 4888 5075
rect 4854 4973 4888 5007
rect 4854 4905 4888 4939
rect 5030 5041 5064 5075
rect 5030 4973 5064 5007
rect 5030 4905 5064 4939
rect 5348 4992 5382 5026
rect 5348 4924 5382 4958
rect 5348 4856 5382 4890
rect 5524 4992 5558 5026
rect 5524 4924 5558 4958
rect 5524 4856 5558 4890
rect 5648 4992 5682 5026
rect 5648 4924 5682 4958
rect 5648 4856 5682 4890
rect 5824 4992 5858 5026
rect 5824 4924 5858 4958
rect 5824 4856 5858 4890
rect 6000 4992 6034 5026
rect 6000 4924 6034 4958
rect 6000 4856 6034 4890
rect 6176 4992 6210 5026
rect 6176 4924 6210 4958
rect 6176 4856 6210 4890
rect 3974 4773 4008 4807
rect 3974 4705 4008 4739
rect 3974 4637 4008 4671
rect 4150 4773 4184 4807
rect 4150 4705 4184 4739
rect 4150 4637 4184 4671
rect 4326 4773 4360 4807
rect 4326 4705 4360 4739
rect 4326 4637 4360 4671
rect 4502 4773 4536 4807
rect 4502 4705 4536 4739
rect 4502 4637 4536 4671
rect 4678 4773 4712 4807
rect 4678 4705 4712 4739
rect 4678 4637 4712 4671
rect 4854 4773 4888 4807
rect 4854 4705 4888 4739
rect 4854 4637 4888 4671
rect 5030 4773 5064 4807
rect 5030 4705 5064 4739
rect 5030 4637 5064 4671
rect 5348 4730 5382 4764
rect 5348 4662 5382 4696
rect 5348 4594 5382 4628
rect 5524 4730 5558 4764
rect 5524 4662 5558 4696
rect 5524 4594 5558 4628
rect 5648 4730 5682 4764
rect 5648 4662 5682 4696
rect 5648 4594 5682 4628
rect 5824 4730 5858 4764
rect 5824 4662 5858 4696
rect 5824 4594 5858 4628
rect 6000 4730 6034 4764
rect 6000 4662 6034 4696
rect 6000 4594 6034 4628
rect 6176 4730 6210 4764
rect 6176 4662 6210 4696
rect 6176 4594 6210 4628
rect 5323 4340 5357 4374
rect 3941 4232 3975 4266
rect 3941 4164 3975 4198
rect 3941 4096 3975 4130
rect 4117 4232 4151 4266
rect 4117 4164 4151 4198
rect 4117 4096 4151 4130
rect 4293 4232 4327 4266
rect 4293 4164 4327 4198
rect 4293 4096 4327 4130
rect 4469 4232 4503 4266
rect 4469 4164 4503 4198
rect 4469 4096 4503 4130
rect 4645 4232 4679 4266
rect 4645 4164 4679 4198
rect 4645 4096 4679 4130
rect 4821 4232 4855 4266
rect 4821 4164 4855 4198
rect 4821 4096 4855 4130
rect 4997 4232 5031 4266
rect 4997 4164 5031 4198
rect 5323 4272 5357 4306
rect 5323 4204 5357 4238
rect 5499 4340 5533 4374
rect 5499 4272 5533 4306
rect 5499 4204 5533 4238
rect 5675 4340 5709 4374
rect 5675 4272 5709 4306
rect 5675 4204 5709 4238
rect 5851 4340 5885 4374
rect 5851 4272 5885 4306
rect 5851 4204 5885 4238
rect 6027 4340 6061 4374
rect 6027 4272 6061 4306
rect 6027 4204 6061 4238
rect 6203 4340 6237 4374
rect 6203 4272 6237 4306
rect 6203 4204 6237 4238
rect 4997 4096 5031 4130
rect 5323 4078 5357 4112
rect 3941 3964 3975 3998
rect 3941 3896 3975 3930
rect 3941 3828 3975 3862
rect 4117 3964 4151 3998
rect 4117 3896 4151 3930
rect 4117 3828 4151 3862
rect 4293 3964 4327 3998
rect 4293 3896 4327 3930
rect 4293 3828 4327 3862
rect 4469 3964 4503 3998
rect 4469 3896 4503 3930
rect 4469 3828 4503 3862
rect 4645 3964 4679 3998
rect 4645 3896 4679 3930
rect 4645 3828 4679 3862
rect 4821 3964 4855 3998
rect 4821 3896 4855 3930
rect 4821 3828 4855 3862
rect 4997 3964 5031 3998
rect 4997 3896 5031 3930
rect 5323 4010 5357 4044
rect 5323 3942 5357 3976
rect 5499 4078 5533 4112
rect 5499 4010 5533 4044
rect 5675 4078 5709 4112
rect 5675 4010 5709 4044
rect 5675 3942 5709 3976
rect 5851 4078 5885 4112
rect 5851 4010 5885 4044
rect 5851 3942 5885 3976
rect 6027 4078 6061 4112
rect 6027 4010 6061 4044
rect 6027 3942 6061 3976
rect 6203 4078 6237 4112
rect 6203 4010 6237 4044
rect 6203 3942 6237 3976
rect 4997 3828 5031 3862
rect -9272 2800 -9238 2834
rect -9272 2732 -9238 2766
rect -9272 2664 -9238 2698
rect -9096 2800 -9062 2834
rect -9096 2732 -9062 2766
rect -9096 2664 -9062 2698
rect -8920 2800 -8886 2834
rect -8920 2732 -8886 2766
rect -8920 2664 -8886 2698
rect -8744 2800 -8710 2834
rect -8744 2732 -8710 2766
rect -8744 2664 -8710 2698
rect -8568 2800 -8534 2834
rect -8568 2732 -8534 2766
rect -8568 2664 -8534 2698
rect -9272 2538 -9238 2572
rect -9272 2470 -9238 2504
rect -9272 2402 -9238 2436
rect -9096 2538 -9062 2572
rect -9096 2470 -9062 2504
rect -8920 2538 -8886 2572
rect -8920 2470 -8886 2504
rect -8920 2402 -8886 2436
rect -8744 2538 -8710 2572
rect -8744 2470 -8710 2504
rect -8744 2402 -8710 2436
rect -8568 2538 -8534 2572
rect -8568 2470 -8534 2504
rect -8568 2402 -8534 2436
<< mvpsubdiff >>
rect 3871 7582 3895 7616
rect 3929 7582 3963 7616
rect 3997 7582 4031 7616
rect 4065 7582 4099 7616
rect 4133 7582 4167 7616
rect 4201 7582 4235 7616
rect 4269 7582 4303 7616
rect 4337 7582 4371 7616
rect 4405 7582 4439 7616
rect 4473 7582 4507 7616
rect 4541 7582 4575 7616
rect 4609 7582 4643 7616
rect 4677 7582 4711 7616
rect 4745 7582 4779 7616
rect 4813 7582 4847 7616
rect 4881 7582 4915 7616
rect 4949 7582 4983 7616
rect 5017 7582 5051 7616
rect 5085 7582 5119 7616
rect 5153 7582 5187 7616
rect 5221 7582 5255 7616
rect 5289 7582 5323 7616
rect 5357 7582 5391 7616
rect 5425 7582 5459 7616
rect 5493 7582 5527 7616
rect 5561 7582 5595 7616
rect 5629 7582 5663 7616
rect 5697 7582 5731 7616
rect 5765 7582 5799 7616
rect 5833 7582 5867 7616
rect 5901 7582 5935 7616
rect 5969 7582 6003 7616
rect 6037 7582 6071 7616
rect 6105 7582 6139 7616
rect 6173 7582 6233 7616
rect 3868 5620 3892 5654
rect 3926 5620 3960 5654
rect 3994 5620 4028 5654
rect 4062 5620 4096 5654
rect 4130 5620 4164 5654
rect 4198 5620 4232 5654
rect 4266 5620 4300 5654
rect 4334 5620 4368 5654
rect 4402 5620 4436 5654
rect 4470 5620 4504 5654
rect 4538 5620 4572 5654
rect 4606 5620 4640 5654
rect 4674 5620 4708 5654
rect 4742 5620 4776 5654
rect 4810 5620 4844 5654
rect 4878 5620 4912 5654
rect 4946 5620 4980 5654
rect 5014 5620 5048 5654
rect 5082 5620 5116 5654
rect 5150 5620 5184 5654
rect 5218 5620 5252 5654
rect 5286 5620 5320 5654
rect 5354 5620 5388 5654
rect 5422 5620 5456 5654
rect 5490 5620 5524 5654
rect 5558 5620 5592 5654
rect 5626 5620 5660 5654
rect 5694 5620 5728 5654
rect 5762 5620 5796 5654
rect 5830 5620 5864 5654
rect 5898 5620 5932 5654
rect 5966 5620 6000 5654
rect 6034 5620 6068 5654
rect 6102 5620 6136 5654
rect 6170 5620 6254 5654
rect 5324 5581 6254 5620
rect 5324 5547 5348 5581
rect 5382 5547 5416 5581
rect 5450 5547 5484 5581
rect 5518 5547 5552 5581
rect 5586 5547 5620 5581
rect 5654 5547 5688 5581
rect 5722 5547 5756 5581
rect 5790 5547 5824 5581
rect 5858 5547 5892 5581
rect 5926 5547 5960 5581
rect 5994 5547 6028 5581
rect 6062 5547 6096 5581
rect 6130 5547 6164 5581
rect 6198 5547 6254 5581
rect 5324 5507 6254 5547
rect 5324 5473 5348 5507
rect 5382 5473 5416 5507
rect 5450 5473 5484 5507
rect 5518 5473 5552 5507
rect 5586 5473 5620 5507
rect 5654 5473 5688 5507
rect 5722 5473 5756 5507
rect 5790 5473 5824 5507
rect 5858 5473 5892 5507
rect 5926 5473 5960 5507
rect 5994 5473 6028 5507
rect 6062 5473 6096 5507
rect 6130 5473 6164 5507
rect 6198 5473 6254 5507
rect 5114 3478 5138 3512
rect 5172 3478 5206 3512
rect 5240 3478 5274 3512
rect 5308 3478 5342 3512
rect 5376 3478 5410 3512
rect 5444 3478 5478 3512
rect 5512 3478 5546 3512
rect 5580 3478 5614 3512
rect 5648 3478 5682 3512
rect 5716 3478 5750 3512
rect 5784 3478 5818 3512
rect 5852 3478 5886 3512
rect 5920 3478 5954 3512
rect 5988 3478 6022 3512
rect 6056 3478 6090 3512
rect 6124 3478 6158 3512
rect 6192 3478 6265 3512
rect 5114 3444 5148 3478
rect 5114 3384 5148 3410
<< mvnsubdiff >>
rect 3871 6601 3895 6635
rect 3929 6601 3963 6635
rect 3997 6601 4031 6635
rect 4065 6601 4099 6635
rect 4133 6601 4167 6635
rect 4201 6601 4235 6635
rect 4269 6601 4303 6635
rect 4337 6601 4371 6635
rect 4405 6601 4439 6635
rect 4473 6601 4507 6635
rect 4541 6601 4575 6635
rect 4609 6601 4643 6635
rect 4677 6601 4711 6635
rect 4745 6601 4779 6635
rect 4813 6601 4847 6635
rect 4881 6601 4915 6635
rect 4949 6601 4983 6635
rect 5017 6601 5051 6635
rect 5085 6601 5119 6635
rect 5153 6601 5187 6635
rect 5221 6601 5255 6635
rect 5289 6601 5323 6635
rect 5357 6601 5391 6635
rect 5425 6601 5459 6635
rect 5493 6601 5527 6635
rect 5561 6601 5595 6635
rect 5629 6601 5663 6635
rect 5697 6601 5731 6635
rect 5765 6601 5799 6635
rect 5833 6601 5867 6635
rect 5901 6601 5935 6635
rect 5969 6601 6003 6635
rect 6037 6601 6071 6635
rect 6105 6601 6139 6635
rect 6173 6601 6229 6635
rect 5194 4470 5230 4501
rect 3996 4436 4035 4470
rect 4069 4436 4103 4470
rect 4137 4436 4171 4470
rect 4205 4436 4239 4470
rect 4273 4436 4307 4470
rect 4341 4436 4375 4470
rect 4409 4436 4443 4470
rect 4477 4436 4511 4470
rect 4545 4436 4579 4470
rect 4613 4436 4647 4470
rect 4681 4436 4715 4470
rect 4749 4436 4783 4470
rect 4817 4436 4851 4470
rect 4885 4436 4919 4470
rect 4953 4436 4987 4470
rect 5021 4436 5055 4470
rect 5089 4436 5123 4470
rect 5157 4467 5230 4470
rect 5264 4467 5298 4501
rect 5332 4467 5366 4501
rect 5400 4467 5434 4501
rect 5468 4467 5502 4501
rect 5536 4467 5570 4501
rect 5604 4467 5638 4501
rect 5672 4467 5706 4501
rect 5740 4467 5774 4501
rect 5808 4467 5842 4501
rect 5876 4467 5910 4501
rect 5944 4467 5978 4501
rect 6012 4467 6046 4501
rect 6080 4467 6114 4501
rect 6148 4467 6218 4501
rect 5157 4436 5228 4467
<< mvpsubdiffcont >>
rect 3895 7582 3929 7616
rect 3963 7582 3997 7616
rect 4031 7582 4065 7616
rect 4099 7582 4133 7616
rect 4167 7582 4201 7616
rect 4235 7582 4269 7616
rect 4303 7582 4337 7616
rect 4371 7582 4405 7616
rect 4439 7582 4473 7616
rect 4507 7582 4541 7616
rect 4575 7582 4609 7616
rect 4643 7582 4677 7616
rect 4711 7582 4745 7616
rect 4779 7582 4813 7616
rect 4847 7582 4881 7616
rect 4915 7582 4949 7616
rect 4983 7582 5017 7616
rect 5051 7582 5085 7616
rect 5119 7582 5153 7616
rect 5187 7582 5221 7616
rect 5255 7582 5289 7616
rect 5323 7582 5357 7616
rect 5391 7582 5425 7616
rect 5459 7582 5493 7616
rect 5527 7582 5561 7616
rect 5595 7582 5629 7616
rect 5663 7582 5697 7616
rect 5731 7582 5765 7616
rect 5799 7582 5833 7616
rect 5867 7582 5901 7616
rect 5935 7582 5969 7616
rect 6003 7582 6037 7616
rect 6071 7582 6105 7616
rect 6139 7582 6173 7616
rect 3892 5620 3926 5654
rect 3960 5620 3994 5654
rect 4028 5620 4062 5654
rect 4096 5620 4130 5654
rect 4164 5620 4198 5654
rect 4232 5620 4266 5654
rect 4300 5620 4334 5654
rect 4368 5620 4402 5654
rect 4436 5620 4470 5654
rect 4504 5620 4538 5654
rect 4572 5620 4606 5654
rect 4640 5620 4674 5654
rect 4708 5620 4742 5654
rect 4776 5620 4810 5654
rect 4844 5620 4878 5654
rect 4912 5620 4946 5654
rect 4980 5620 5014 5654
rect 5048 5620 5082 5654
rect 5116 5620 5150 5654
rect 5184 5620 5218 5654
rect 5252 5620 5286 5654
rect 5320 5620 5354 5654
rect 5388 5620 5422 5654
rect 5456 5620 5490 5654
rect 5524 5620 5558 5654
rect 5592 5620 5626 5654
rect 5660 5620 5694 5654
rect 5728 5620 5762 5654
rect 5796 5620 5830 5654
rect 5864 5620 5898 5654
rect 5932 5620 5966 5654
rect 6000 5620 6034 5654
rect 6068 5620 6102 5654
rect 6136 5620 6170 5654
rect 5348 5547 5382 5581
rect 5416 5547 5450 5581
rect 5484 5547 5518 5581
rect 5552 5547 5586 5581
rect 5620 5547 5654 5581
rect 5688 5547 5722 5581
rect 5756 5547 5790 5581
rect 5824 5547 5858 5581
rect 5892 5547 5926 5581
rect 5960 5547 5994 5581
rect 6028 5547 6062 5581
rect 6096 5547 6130 5581
rect 6164 5547 6198 5581
rect 5348 5473 5382 5507
rect 5416 5473 5450 5507
rect 5484 5473 5518 5507
rect 5552 5473 5586 5507
rect 5620 5473 5654 5507
rect 5688 5473 5722 5507
rect 5756 5473 5790 5507
rect 5824 5473 5858 5507
rect 5892 5473 5926 5507
rect 5960 5473 5994 5507
rect 6028 5473 6062 5507
rect 6096 5473 6130 5507
rect 6164 5473 6198 5507
rect 5138 3478 5172 3512
rect 5206 3478 5240 3512
rect 5274 3478 5308 3512
rect 5342 3478 5376 3512
rect 5410 3478 5444 3512
rect 5478 3478 5512 3512
rect 5546 3478 5580 3512
rect 5614 3478 5648 3512
rect 5682 3478 5716 3512
rect 5750 3478 5784 3512
rect 5818 3478 5852 3512
rect 5886 3478 5920 3512
rect 5954 3478 5988 3512
rect 6022 3478 6056 3512
rect 6090 3478 6124 3512
rect 6158 3478 6192 3512
rect 5114 3410 5148 3444
<< mvnsubdiffcont >>
rect 3895 6601 3929 6635
rect 3963 6601 3997 6635
rect 4031 6601 4065 6635
rect 4099 6601 4133 6635
rect 4167 6601 4201 6635
rect 4235 6601 4269 6635
rect 4303 6601 4337 6635
rect 4371 6601 4405 6635
rect 4439 6601 4473 6635
rect 4507 6601 4541 6635
rect 4575 6601 4609 6635
rect 4643 6601 4677 6635
rect 4711 6601 4745 6635
rect 4779 6601 4813 6635
rect 4847 6601 4881 6635
rect 4915 6601 4949 6635
rect 4983 6601 5017 6635
rect 5051 6601 5085 6635
rect 5119 6601 5153 6635
rect 5187 6601 5221 6635
rect 5255 6601 5289 6635
rect 5323 6601 5357 6635
rect 5391 6601 5425 6635
rect 5459 6601 5493 6635
rect 5527 6601 5561 6635
rect 5595 6601 5629 6635
rect 5663 6601 5697 6635
rect 5731 6601 5765 6635
rect 5799 6601 5833 6635
rect 5867 6601 5901 6635
rect 5935 6601 5969 6635
rect 6003 6601 6037 6635
rect 6071 6601 6105 6635
rect 6139 6601 6173 6635
rect 4035 4436 4069 4470
rect 4103 4436 4137 4470
rect 4171 4436 4205 4470
rect 4239 4436 4273 4470
rect 4307 4436 4341 4470
rect 4375 4436 4409 4470
rect 4443 4436 4477 4470
rect 4511 4436 4545 4470
rect 4579 4436 4613 4470
rect 4647 4436 4681 4470
rect 4715 4436 4749 4470
rect 4783 4436 4817 4470
rect 4851 4436 4885 4470
rect 4919 4436 4953 4470
rect 4987 4436 5021 4470
rect 5055 4436 5089 4470
rect 5123 4436 5157 4470
rect 5230 4467 5264 4501
rect 5298 4467 5332 4501
rect 5366 4467 5400 4501
rect 5434 4467 5468 4501
rect 5502 4467 5536 4501
rect 5570 4467 5604 4501
rect 5638 4467 5672 4501
rect 5706 4467 5740 4501
rect 5774 4467 5808 4501
rect 5842 4467 5876 4501
rect 5910 4467 5944 4501
rect 5978 4467 6012 4501
rect 6046 4467 6080 4501
rect 6114 4467 6148 4501
<< poly >>
rect 3924 7508 4044 7534
rect 4100 7508 4220 7534
rect 4400 7508 4520 7534
rect 4576 7508 4696 7534
rect 4752 7508 4872 7534
rect 4928 7508 5048 7534
rect 5228 7508 5348 7534
rect 5404 7508 5524 7534
rect 5704 7508 5824 7534
rect 5880 7508 6000 7534
rect 6056 7508 6176 7534
rect 3924 7320 4044 7368
rect 3924 7286 3969 7320
rect 4003 7286 4044 7320
rect 3924 7252 4044 7286
rect 3924 7218 3969 7252
rect 4003 7218 4044 7252
rect 3924 7170 4044 7218
rect 4100 7320 4220 7368
rect 4100 7286 4140 7320
rect 4174 7286 4220 7320
rect 4100 7252 4220 7286
rect 4100 7218 4140 7252
rect 4174 7218 4220 7252
rect 4100 7170 4220 7218
rect 4400 7320 4520 7368
rect 4400 7286 4445 7320
rect 4479 7286 4520 7320
rect 4400 7252 4520 7286
rect 4400 7218 4445 7252
rect 4479 7218 4520 7252
rect 4400 7170 4520 7218
rect 4576 7320 4696 7368
rect 4576 7286 4616 7320
rect 4650 7286 4696 7320
rect 4576 7252 4696 7286
rect 4576 7218 4616 7252
rect 4650 7218 4696 7252
rect 4576 7170 4696 7218
rect 4752 7320 4872 7368
rect 4752 7286 4798 7320
rect 4832 7286 4872 7320
rect 4752 7252 4872 7286
rect 4752 7218 4798 7252
rect 4832 7218 4872 7252
rect 4752 7170 4872 7218
rect 4928 7320 5048 7368
rect 4928 7286 4969 7320
rect 5003 7286 5048 7320
rect 4928 7252 5048 7286
rect 4928 7218 4969 7252
rect 5003 7218 5048 7252
rect 4928 7170 5048 7218
rect 5228 7320 5348 7368
rect 5228 7286 5273 7320
rect 5307 7286 5348 7320
rect 5228 7252 5348 7286
rect 5228 7218 5273 7252
rect 5307 7218 5348 7252
rect 5228 7170 5348 7218
rect 5404 7320 5524 7368
rect 5404 7286 5444 7320
rect 5478 7286 5524 7320
rect 5404 7252 5524 7286
rect 5404 7218 5444 7252
rect 5478 7218 5524 7252
rect 5404 7170 5524 7218
rect 5704 7320 5824 7368
rect 5704 7286 5746 7320
rect 5780 7286 5824 7320
rect 5704 7252 5824 7286
rect 5704 7218 5746 7252
rect 5780 7218 5824 7252
rect 5704 7170 5824 7218
rect 5880 7342 6000 7368
rect 6056 7342 6176 7368
rect 5880 7320 6176 7342
rect 5880 7286 5918 7320
rect 5952 7286 6105 7320
rect 6139 7286 6176 7320
rect 5880 7252 6176 7286
rect 5880 7218 5918 7252
rect 5952 7218 6105 7252
rect 6139 7218 6176 7252
rect 5880 7196 6176 7218
rect 5880 7170 6000 7196
rect 6056 7170 6176 7196
rect 3924 6902 4044 6970
rect 4100 6902 4220 6970
rect 4400 6902 4520 6970
rect 4576 6902 4696 6970
rect 4752 6902 4872 6970
rect 4928 6902 5048 6970
rect 5228 6902 5348 6970
rect 5404 6902 5524 6970
rect 5704 6902 5824 6970
rect 5880 6902 6000 6970
rect 6056 6902 6176 6970
rect 3924 6676 4044 6702
rect 4100 6676 4220 6702
rect 4400 6676 4520 6702
rect 4576 6676 4696 6702
rect 4752 6676 4872 6702
rect 4928 6676 5048 6702
rect 5228 6676 5348 6702
rect 5404 6676 5524 6702
rect 5704 6676 5824 6702
rect 5880 6676 6000 6702
rect 6056 6676 6176 6702
rect 3924 6534 4044 6560
rect 4100 6534 4220 6560
rect 4400 6534 4520 6560
rect 4576 6534 4696 6560
rect 4876 6534 4996 6560
rect 5052 6534 5172 6560
rect 5228 6534 5348 6560
rect 5404 6534 5524 6560
rect 5704 6534 5824 6560
rect 5880 6534 6000 6560
rect 6056 6534 6176 6560
rect 3924 6266 4044 6334
rect 4100 6266 4220 6334
rect 4400 6266 4520 6334
rect 4576 6266 4696 6334
rect 4876 6266 4996 6334
rect 5052 6266 5172 6334
rect 5228 6266 5348 6334
rect 5404 6266 5524 6334
rect 5704 6266 5824 6334
rect 5880 6266 6000 6334
rect 6056 6266 6176 6334
rect 3924 6018 4044 6066
rect 3924 5984 3965 6018
rect 3999 5984 4044 6018
rect 3924 5950 4044 5984
rect 3924 5916 3965 5950
rect 3999 5916 4044 5950
rect 3924 5868 4044 5916
rect 4100 6018 4220 6066
rect 4100 5984 4143 6018
rect 4177 5984 4220 6018
rect 4100 5950 4220 5984
rect 4100 5916 4143 5950
rect 4177 5916 4220 5950
rect 4100 5868 4220 5916
rect 4400 6018 4520 6066
rect 4400 5984 4446 6018
rect 4480 5984 4520 6018
rect 4400 5950 4520 5984
rect 4400 5916 4446 5950
rect 4480 5916 4520 5950
rect 4400 5868 4520 5916
rect 4576 6018 4696 6066
rect 4576 5984 4617 6018
rect 4651 5984 4696 6018
rect 4576 5950 4696 5984
rect 4576 5916 4617 5950
rect 4651 5916 4696 5950
rect 4576 5868 4696 5916
rect 4876 6018 4996 6066
rect 4876 5984 4921 6018
rect 4955 5984 4996 6018
rect 4876 5950 4996 5984
rect 4876 5916 4921 5950
rect 4955 5916 4996 5950
rect 4876 5868 4996 5916
rect 5052 6018 5172 6066
rect 5052 5984 5092 6018
rect 5126 5984 5172 6018
rect 5052 5950 5172 5984
rect 5052 5916 5092 5950
rect 5126 5916 5172 5950
rect 5052 5868 5172 5916
rect 5228 6018 5348 6066
rect 5228 5984 5274 6018
rect 5308 5984 5348 6018
rect 5228 5950 5348 5984
rect 5228 5916 5274 5950
rect 5308 5916 5348 5950
rect 5228 5868 5348 5916
rect 5404 6018 5524 6066
rect 5404 5984 5445 6018
rect 5479 5984 5524 6018
rect 5404 5950 5524 5984
rect 5404 5916 5445 5950
rect 5479 5916 5524 5950
rect 5404 5868 5524 5916
rect 5704 6018 5824 6066
rect 5704 5984 5746 6018
rect 5780 5984 5824 6018
rect 5704 5950 5824 5984
rect 5704 5916 5746 5950
rect 5780 5916 5824 5950
rect 5704 5868 5824 5916
rect 5880 6040 6000 6066
rect 6056 6040 6176 6066
rect 5880 6018 6176 6040
rect 5880 5984 5917 6018
rect 5951 5984 6104 6018
rect 6138 5984 6176 6018
rect 5880 5950 6176 5984
rect 5880 5916 5917 5950
rect 5951 5916 6104 5950
rect 6138 5916 6176 5950
rect 5880 5894 6176 5916
rect 5880 5868 6000 5894
rect 6056 5868 6176 5894
rect 3924 5702 4044 5728
rect 4100 5702 4220 5728
rect 4400 5702 4520 5728
rect 4576 5702 4696 5728
rect 4876 5702 4996 5728
rect 5052 5702 5172 5728
rect 5228 5702 5348 5728
rect 5404 5702 5524 5728
rect 5704 5702 5824 5728
rect 5880 5702 6000 5728
rect 6056 5702 6176 5728
rect 4019 5565 4315 5581
rect 4019 5531 4035 5565
rect 4069 5531 4112 5565
rect 4146 5531 4189 5565
rect 4223 5531 4265 5565
rect 4299 5531 4315 5565
rect 4019 5515 4315 5531
rect 4363 5565 4497 5581
rect 4363 5531 4379 5565
rect 4413 5531 4447 5565
rect 4481 5531 4497 5565
rect 4363 5515 4497 5531
rect 4891 5565 5025 5581
rect 4891 5531 4907 5565
rect 4941 5531 4975 5565
rect 5009 5531 5025 5565
rect 4891 5515 5025 5531
rect 4019 5489 4139 5515
rect 4195 5489 4315 5515
rect 4371 5489 4491 5515
rect 4547 5489 4667 5515
rect 4723 5489 4843 5515
rect 4899 5489 5019 5515
rect 5393 5382 5513 5408
rect 5693 5382 5813 5408
rect 5869 5382 5989 5408
rect 6045 5382 6165 5408
rect 4019 5087 4139 5349
rect 4195 5087 4315 5349
rect 4371 5323 4491 5349
rect 4547 5281 4667 5349
rect 4371 5247 4667 5281
rect 4371 5213 4413 5247
rect 4447 5242 4667 5247
rect 4447 5213 4491 5242
rect 4371 5179 4491 5213
rect 4723 5200 4843 5349
rect 4371 5145 4413 5179
rect 4447 5145 4491 5179
rect 4371 5087 4491 5145
rect 4547 5161 4843 5200
rect 4547 5087 4667 5161
rect 4723 5087 4843 5119
rect 4899 5087 5019 5349
rect 5393 5194 5513 5242
rect 5393 5160 5437 5194
rect 5471 5160 5513 5194
rect 5393 5126 5513 5160
rect 5393 5092 5437 5126
rect 5471 5092 5513 5126
rect 5393 5044 5513 5092
rect 5693 5216 5813 5242
rect 5869 5216 5989 5242
rect 5693 5194 5989 5216
rect 5693 5160 5731 5194
rect 5765 5160 5918 5194
rect 5952 5160 5989 5194
rect 5693 5126 5989 5160
rect 5693 5092 5731 5126
rect 5765 5092 5918 5126
rect 5952 5092 5989 5126
rect 5693 5070 5989 5092
rect 5693 5044 5813 5070
rect 5869 5044 5989 5070
rect 6045 5194 6165 5242
rect 6045 5160 6089 5194
rect 6123 5160 6165 5194
rect 6045 5126 6165 5160
rect 6045 5092 6089 5126
rect 6123 5092 6165 5126
rect 6045 5044 6165 5092
rect 4019 4819 4139 4887
rect 4195 4819 4315 4887
rect 4371 4819 4491 4887
rect 4547 4819 4667 4887
rect 4723 4819 4843 4887
rect 4899 4819 5019 4887
rect 5393 4776 5513 4844
rect 5693 4776 5813 4844
rect 5869 4776 5989 4844
rect 6045 4776 6165 4844
rect 4019 4587 4139 4619
rect 4195 4587 4315 4619
rect 4371 4587 4491 4619
rect 4547 4587 4667 4619
rect 4723 4587 4843 4619
rect 4899 4587 5019 4619
rect 4019 4571 4315 4587
rect 4019 4537 4035 4571
rect 4069 4537 4112 4571
rect 4146 4537 4189 4571
rect 4223 4537 4265 4571
rect 4299 4537 4315 4571
rect 4019 4521 4315 4537
rect 4539 4571 4673 4587
rect 4539 4537 4555 4571
rect 4589 4537 4623 4571
rect 4657 4537 4673 4571
rect 4539 4521 4673 4537
rect 4723 4571 5019 4587
rect 4723 4537 4739 4571
rect 4773 4537 4816 4571
rect 4850 4537 4893 4571
rect 4927 4537 4969 4571
rect 5003 4537 5019 4571
rect 5393 4550 5513 4576
rect 5693 4550 5813 4576
rect 5869 4550 5989 4576
rect 6045 4550 6165 4576
rect 4723 4521 5019 4537
rect 5368 4392 5488 4418
rect 5544 4392 5664 4418
rect 5720 4392 5840 4418
rect 5896 4392 6016 4418
rect 6072 4392 6192 4418
rect 3986 4366 4282 4382
rect 3986 4332 4002 4366
rect 4036 4332 4079 4366
rect 4113 4332 4156 4366
rect 4190 4332 4232 4366
rect 4266 4332 4282 4366
rect 3986 4316 4282 4332
rect 4506 4366 4640 4382
rect 4506 4332 4522 4366
rect 4556 4332 4590 4366
rect 4624 4332 4640 4366
rect 4506 4316 4640 4332
rect 4690 4366 4986 4382
rect 4690 4332 4706 4366
rect 4740 4332 4783 4366
rect 4817 4332 4860 4366
rect 4894 4332 4936 4366
rect 4970 4332 4986 4366
rect 4690 4316 4986 4332
rect 3986 4284 4106 4316
rect 4162 4284 4282 4316
rect 4338 4284 4458 4316
rect 4514 4284 4634 4316
rect 4690 4284 4810 4316
rect 4866 4284 4986 4316
rect 5368 4124 5488 4192
rect 5544 4124 5664 4192
rect 5720 4124 5840 4192
rect 5896 4124 6016 4192
rect 6072 4124 6192 4192
rect 3986 4016 4106 4084
rect 4162 4016 4282 4084
rect 4338 4016 4458 4084
rect 4514 4016 4634 4084
rect 4690 4016 4810 4084
rect 4866 4016 4986 4084
rect 5368 3876 5488 3924
rect 5368 3842 5409 3876
rect 5443 3842 5488 3876
rect 3986 3554 4106 3816
rect 4162 3554 4282 3816
rect 4338 3758 4458 3816
rect 4338 3724 4380 3758
rect 4414 3724 4458 3758
rect 4338 3690 4458 3724
rect 4338 3656 4380 3690
rect 4414 3656 4458 3690
rect 4514 3742 4634 3816
rect 4690 3784 4810 3816
rect 4514 3709 4810 3742
rect 4514 3675 4553 3709
rect 4587 3675 4621 3709
rect 4655 3675 4810 3709
rect 4514 3659 4810 3675
rect 4338 3622 4458 3656
rect 4338 3554 4458 3580
rect 4514 3554 4634 3580
rect 4690 3554 4810 3659
rect 4866 3554 4986 3816
rect 5368 3808 5488 3842
rect 5368 3774 5409 3808
rect 5443 3774 5488 3808
rect 5368 3726 5488 3774
rect 5544 3876 5664 3924
rect 5544 3842 5587 3876
rect 5621 3842 5664 3876
rect 5544 3808 5664 3842
rect 5544 3774 5587 3808
rect 5621 3774 5664 3808
rect 5544 3726 5664 3774
rect 5720 3898 5840 3924
rect 5896 3898 6016 3924
rect 5720 3876 6016 3898
rect 5720 3842 5758 3876
rect 5792 3842 5945 3876
rect 5979 3842 6016 3876
rect 5720 3808 6016 3842
rect 5720 3774 5758 3808
rect 5792 3774 5945 3808
rect 5979 3774 6016 3808
rect 5720 3752 6016 3774
rect 5720 3726 5840 3752
rect 5896 3726 6016 3752
rect 6072 3876 6192 3924
rect 6072 3842 6116 3876
rect 6150 3842 6192 3876
rect 6072 3808 6192 3842
rect 6072 3774 6116 3808
rect 6150 3774 6192 3808
rect 6072 3726 6192 3774
rect 5368 3560 5488 3586
rect 5544 3560 5664 3586
rect 5720 3560 5840 3586
rect 5896 3560 6016 3586
rect 6072 3560 6192 3586
rect 3986 3388 4106 3414
rect 4162 3388 4282 3414
rect 4338 3388 4458 3414
rect 4514 3388 4634 3414
rect 4690 3388 4810 3414
rect 4866 3388 4986 3414
rect 3986 3372 4282 3388
rect 3986 3338 4002 3372
rect 4036 3338 4079 3372
rect 4113 3338 4156 3372
rect 4190 3338 4232 3372
rect 4266 3338 4282 3372
rect 3986 3322 4282 3338
rect 4330 3372 4464 3388
rect 4330 3338 4346 3372
rect 4380 3338 4414 3372
rect 4448 3338 4464 3372
rect 4330 3322 4464 3338
rect 4858 3372 4992 3388
rect 4858 3338 4874 3372
rect 4908 3338 4942 3372
rect 4976 3338 4992 3372
rect 4858 3322 4992 3338
rect -9227 2852 -9107 2878
rect -9051 2852 -8931 2878
rect -8875 2852 -8755 2878
rect -8699 2852 -8579 2878
rect -9227 2584 -9107 2652
rect -9051 2584 -8931 2652
rect -8875 2584 -8755 2652
rect -8699 2584 -8579 2652
rect -9227 2336 -9107 2384
rect -9227 2302 -9186 2336
rect -9152 2302 -9107 2336
rect -9227 2268 -9107 2302
rect -9227 2234 -9186 2268
rect -9152 2234 -9107 2268
rect -9227 2186 -9107 2234
rect -9051 2336 -8931 2384
rect -9051 2302 -9008 2336
rect -8974 2302 -8931 2336
rect -9051 2268 -8931 2302
rect -9051 2234 -9008 2268
rect -8974 2234 -8931 2268
rect -9051 2186 -8931 2234
rect -8875 2336 -8755 2384
rect -8875 2302 -8829 2336
rect -8795 2302 -8755 2336
rect -8875 2268 -8755 2302
rect -8875 2234 -8829 2268
rect -8795 2234 -8755 2268
rect -8875 2186 -8755 2234
rect -8699 2336 -8579 2384
rect -8699 2302 -8658 2336
rect -8624 2302 -8579 2336
rect -8699 2268 -8579 2302
rect -8699 2234 -8658 2268
rect -8624 2234 -8579 2268
rect -8699 2186 -8579 2234
rect -9227 2020 -9107 2046
rect -9051 2020 -8931 2046
rect -8875 2020 -8755 2046
rect -8699 2020 -8579 2046
<< polycont >>
rect 3969 7286 4003 7320
rect 3969 7218 4003 7252
rect 4140 7286 4174 7320
rect 4140 7218 4174 7252
rect 4445 7286 4479 7320
rect 4445 7218 4479 7252
rect 4616 7286 4650 7320
rect 4616 7218 4650 7252
rect 4798 7286 4832 7320
rect 4798 7218 4832 7252
rect 4969 7286 5003 7320
rect 4969 7218 5003 7252
rect 5273 7286 5307 7320
rect 5273 7218 5307 7252
rect 5444 7286 5478 7320
rect 5444 7218 5478 7252
rect 5746 7286 5780 7320
rect 5746 7218 5780 7252
rect 5918 7286 5952 7320
rect 6105 7286 6139 7320
rect 5918 7218 5952 7252
rect 6105 7218 6139 7252
rect 3965 5984 3999 6018
rect 3965 5916 3999 5950
rect 4143 5984 4177 6018
rect 4143 5916 4177 5950
rect 4446 5984 4480 6018
rect 4446 5916 4480 5950
rect 4617 5984 4651 6018
rect 4617 5916 4651 5950
rect 4921 5984 4955 6018
rect 4921 5916 4955 5950
rect 5092 5984 5126 6018
rect 5092 5916 5126 5950
rect 5274 5984 5308 6018
rect 5274 5916 5308 5950
rect 5445 5984 5479 6018
rect 5445 5916 5479 5950
rect 5746 5984 5780 6018
rect 5746 5916 5780 5950
rect 5917 5984 5951 6018
rect 6104 5984 6138 6018
rect 5917 5916 5951 5950
rect 6104 5916 6138 5950
rect 4035 5531 4069 5565
rect 4112 5531 4146 5565
rect 4189 5531 4223 5565
rect 4265 5531 4299 5565
rect 4379 5531 4413 5565
rect 4447 5531 4481 5565
rect 4907 5531 4941 5565
rect 4975 5531 5009 5565
rect 4413 5213 4447 5247
rect 4413 5145 4447 5179
rect 5437 5160 5471 5194
rect 5437 5092 5471 5126
rect 5731 5160 5765 5194
rect 5918 5160 5952 5194
rect 5731 5092 5765 5126
rect 5918 5092 5952 5126
rect 6089 5160 6123 5194
rect 6089 5092 6123 5126
rect 4035 4537 4069 4571
rect 4112 4537 4146 4571
rect 4189 4537 4223 4571
rect 4265 4537 4299 4571
rect 4555 4537 4589 4571
rect 4623 4537 4657 4571
rect 4739 4537 4773 4571
rect 4816 4537 4850 4571
rect 4893 4537 4927 4571
rect 4969 4537 5003 4571
rect 4002 4332 4036 4366
rect 4079 4332 4113 4366
rect 4156 4332 4190 4366
rect 4232 4332 4266 4366
rect 4522 4332 4556 4366
rect 4590 4332 4624 4366
rect 4706 4332 4740 4366
rect 4783 4332 4817 4366
rect 4860 4332 4894 4366
rect 4936 4332 4970 4366
rect 5409 3842 5443 3876
rect 4380 3724 4414 3758
rect 4380 3656 4414 3690
rect 4553 3675 4587 3709
rect 4621 3675 4655 3709
rect 5409 3774 5443 3808
rect 5587 3842 5621 3876
rect 5587 3774 5621 3808
rect 5758 3842 5792 3876
rect 5945 3842 5979 3876
rect 5758 3774 5792 3808
rect 5945 3774 5979 3808
rect 6116 3842 6150 3876
rect 6116 3774 6150 3808
rect 4002 3338 4036 3372
rect 4079 3338 4113 3372
rect 4156 3338 4190 3372
rect 4232 3338 4266 3372
rect 4346 3338 4380 3372
rect 4414 3338 4448 3372
rect 4874 3338 4908 3372
rect 4942 3338 4976 3372
rect -9186 2302 -9152 2336
rect -9186 2234 -9152 2268
rect -9008 2302 -8974 2336
rect -9008 2234 -8974 2268
rect -8829 2302 -8795 2336
rect -8829 2234 -8795 2268
rect -8658 2302 -8624 2336
rect -8658 2234 -8624 2268
<< locali >>
rect 3871 7582 3883 7616
rect 3929 7582 3955 7616
rect 3997 7582 4027 7616
rect 4065 7582 4099 7616
rect 4133 7582 4167 7616
rect 4205 7582 4235 7616
rect 4277 7582 4303 7616
rect 4349 7582 4371 7616
rect 4421 7582 4439 7616
rect 4493 7582 4507 7616
rect 4565 7582 4575 7616
rect 4637 7582 4643 7616
rect 4709 7582 4711 7616
rect 4745 7582 4747 7616
rect 4813 7582 4819 7616
rect 4881 7582 4891 7616
rect 4949 7582 4963 7616
rect 5017 7582 5035 7616
rect 5085 7582 5107 7616
rect 5153 7582 5179 7616
rect 5221 7582 5251 7616
rect 5289 7582 5323 7616
rect 5357 7582 5391 7616
rect 5429 7582 5459 7616
rect 5501 7582 5527 7616
rect 5573 7582 5595 7616
rect 5645 7582 5663 7616
rect 5717 7582 5731 7616
rect 5789 7582 5799 7616
rect 5861 7582 5867 7616
rect 5933 7582 5935 7616
rect 5969 7582 5971 7616
rect 6037 7582 6043 7616
rect 6105 7582 6115 7616
rect 6173 7582 6187 7616
rect 6221 7582 6233 7616
rect 3879 7482 3918 7498
rect 3913 7448 3918 7482
rect 3879 7425 3918 7448
rect 4231 7482 4265 7497
rect 3879 7414 4089 7425
rect 3913 7391 4089 7414
rect 3879 7364 3913 7380
rect 3953 7286 3969 7320
rect 4003 7302 4019 7320
rect 3953 7268 3971 7286
rect 4005 7268 4019 7302
rect 3953 7252 4019 7268
rect 3953 7218 3969 7252
rect 4003 7230 4019 7252
rect 4005 7218 4019 7230
rect 3879 7152 3913 7168
rect 3879 7084 3913 7118
rect 3879 7016 3913 7050
rect 3879 6890 3913 6982
rect 3879 6822 3913 6856
rect 3879 6780 3913 6788
rect 3879 6708 3913 6720
rect 4055 7152 4089 7391
rect 4231 7414 4265 7425
rect 4231 7364 4265 7380
rect 4355 7482 4394 7498
rect 4389 7448 4394 7482
rect 4355 7425 4394 7448
rect 4707 7482 4741 7497
rect 5054 7482 5093 7498
rect 5054 7448 5059 7482
rect 5054 7425 5093 7448
rect 4355 7414 4565 7425
rect 4389 7391 4565 7414
rect 4355 7364 4389 7380
rect 4055 7084 4089 7118
rect 4055 7016 4089 7020
rect 4055 6890 4089 6948
rect 4055 6822 4089 6856
rect 4124 7286 4140 7320
rect 4174 7286 4190 7320
rect 4124 7252 4190 7286
rect 4124 7218 4140 7252
rect 4174 7218 4190 7252
rect 4124 6939 4190 7218
rect 4429 7305 4445 7320
rect 4429 7271 4443 7305
rect 4479 7286 4495 7320
rect 4477 7271 4495 7286
rect 4429 7252 4495 7271
rect 4429 7233 4445 7252
rect 4429 7199 4443 7233
rect 4479 7218 4495 7252
rect 4477 7199 4495 7218
rect 4124 6905 4144 6939
rect 4178 6905 4190 6939
rect 4124 6867 4190 6905
rect 4124 6833 4144 6867
rect 4178 6833 4190 6867
rect 4124 6831 4190 6833
rect 4231 7152 4265 7168
rect 4231 7084 4265 7118
rect 4231 7016 4265 7050
rect 4231 6890 4265 6982
rect 4055 6754 4089 6788
rect 4055 6702 4089 6720
rect 4231 6822 4265 6856
rect 4231 6780 4265 6788
rect 4231 6708 4265 6720
rect 4355 7152 4389 7168
rect 4531 7157 4565 7391
rect 4707 7414 4741 7425
rect 4707 7364 4741 7380
rect 4883 7414 5093 7425
rect 4883 7391 5059 7414
rect 4600 7305 4616 7320
rect 4600 7271 4612 7305
rect 4650 7286 4666 7320
rect 4646 7271 4666 7286
rect 4600 7252 4666 7271
rect 4600 7233 4616 7252
rect 4600 7199 4612 7233
rect 4650 7218 4666 7252
rect 4782 7309 4798 7320
rect 4782 7275 4795 7309
rect 4832 7286 4848 7320
rect 4829 7275 4848 7286
rect 4782 7252 4848 7275
rect 4782 7237 4798 7252
rect 4782 7218 4795 7237
rect 4832 7218 4848 7252
rect 4646 7199 4666 7218
rect 4355 7084 4389 7118
rect 4564 7152 4565 7157
rect 4530 7118 4531 7123
rect 4530 7085 4565 7118
rect 4564 7084 4565 7085
rect 4355 7016 4389 7050
rect 4355 6890 4389 6982
rect 4355 6822 4389 6856
rect 4355 6780 4389 6788
rect 4355 6708 4389 6720
rect 4531 7016 4565 7050
rect 4531 6890 4565 6982
rect 4531 6822 4565 6856
rect 4531 6754 4565 6788
rect 4531 6702 4565 6720
rect 4707 7152 4741 7168
rect 4707 7084 4741 7118
rect 4707 7016 4741 7050
rect 4707 6890 4741 6982
rect 4707 6822 4741 6856
rect 4707 6780 4741 6788
rect 4707 6708 4741 6720
rect 4883 7152 4917 7391
rect 5059 7364 5093 7380
rect 5183 7482 5222 7498
rect 5217 7448 5222 7482
rect 5183 7425 5222 7448
rect 5535 7482 5569 7497
rect 5183 7414 5393 7425
rect 5217 7391 5393 7414
rect 5183 7364 5217 7380
rect 4953 7309 4969 7320
rect 4953 7275 4968 7309
rect 5003 7286 5019 7320
rect 5002 7275 5019 7286
rect 4953 7252 5019 7275
rect 4953 7237 4969 7252
rect 4953 7218 4968 7237
rect 5003 7218 5019 7252
rect 5257 7286 5273 7320
rect 5307 7286 5323 7320
rect 5257 7252 5323 7286
rect 5257 7218 5273 7252
rect 5307 7218 5323 7252
rect 4883 7084 4917 7118
rect 4883 7025 4917 7050
rect 4883 6953 4917 6982
rect 4883 6890 4917 6919
rect 4883 6822 4917 6856
rect 4883 6754 4917 6788
rect 4883 6702 4917 6720
rect 5059 7152 5093 7168
rect 5059 7084 5093 7118
rect 5059 7016 5093 7050
rect 5059 6890 5093 6982
rect 5059 6822 5093 6856
rect 5059 6780 5093 6788
rect 5059 6708 5093 6720
rect 5183 7152 5217 7168
rect 5183 7084 5217 7118
rect 5183 7016 5217 7050
rect 5183 6890 5217 6982
rect 5257 7025 5323 7218
rect 5257 6991 5267 7025
rect 5301 6991 5323 7025
rect 5257 6953 5323 6991
rect 5257 6921 5267 6953
rect 5301 6921 5323 6953
rect 5359 7152 5393 7391
rect 5535 7414 5569 7425
rect 5535 7364 5569 7380
rect 5659 7482 5693 7498
rect 5659 7414 5693 7448
rect 5428 7286 5444 7320
rect 5478 7309 5494 7320
rect 5428 7275 5445 7286
rect 5479 7275 5494 7309
rect 5428 7252 5494 7275
rect 5428 7218 5444 7252
rect 5478 7237 5494 7252
rect 5479 7218 5494 7237
rect 5359 7084 5393 7118
rect 5359 7027 5393 7050
rect 5359 6955 5393 6982
rect 5183 6822 5217 6856
rect 5183 6780 5217 6788
rect 5183 6708 5217 6720
rect 5359 6890 5393 6921
rect 5359 6822 5393 6856
rect 5359 6754 5393 6788
rect 5359 6702 5393 6720
rect 5535 7152 5569 7168
rect 5535 7084 5569 7118
rect 5535 7016 5569 7050
rect 5535 6890 5569 6982
rect 5535 6822 5569 6856
rect 5535 6780 5569 6788
rect 5535 6708 5569 6720
rect 5659 7167 5693 7380
rect 5835 7482 5869 7497
rect 5835 7414 5869 7425
rect 5835 7364 5869 7380
rect 6011 7482 6045 7498
rect 6011 7414 6045 7448
rect 5659 7095 5693 7118
rect 5659 7016 5693 7050
rect 5659 6890 5693 6982
rect 5730 7286 5746 7320
rect 5780 7286 5796 7320
rect 5730 7252 5796 7286
rect 5730 7218 5746 7252
rect 5780 7218 5796 7252
rect 5902 7286 5918 7320
rect 5952 7286 5968 7320
rect 5902 7252 5968 7286
rect 5902 7218 5918 7252
rect 5952 7218 5968 7252
rect 5730 7034 5796 7218
rect 5730 7000 5743 7034
rect 5777 7000 5796 7034
rect 5730 6962 5796 7000
rect 5730 6928 5743 6962
rect 5777 6928 5796 6962
rect 5835 7152 5869 7168
rect 5835 7084 5869 7118
rect 5835 7016 5869 7050
rect 5904 7167 5968 7218
rect 5904 7133 5917 7167
rect 5951 7133 5968 7167
rect 5904 7095 5968 7133
rect 5904 7061 5917 7095
rect 5951 7061 5968 7095
rect 5904 7043 5968 7061
rect 6011 7152 6045 7380
rect 6187 7482 6221 7497
rect 6187 7414 6221 7425
rect 6187 7364 6221 7380
rect 6011 7084 6045 7118
rect 5659 6822 5693 6856
rect 5659 6754 5693 6788
rect 5659 6702 5693 6720
rect 5835 6890 5869 6982
rect 5835 6822 5869 6856
rect 5835 6780 5869 6788
rect 5835 6708 5869 6720
rect 6011 7016 6045 7050
rect 6089 7286 6105 7320
rect 6139 7286 6155 7320
rect 6089 7252 6155 7286
rect 6089 7218 6105 7252
rect 6139 7218 6155 7252
rect 6089 7167 6151 7218
rect 6089 7133 6111 7167
rect 6145 7133 6151 7167
rect 6089 7095 6151 7133
rect 6089 7061 6111 7095
rect 6145 7061 6151 7095
rect 6089 7043 6151 7061
rect 6187 7152 6221 7168
rect 6187 7084 6221 7118
rect 6011 6910 6045 6948
rect 6011 6822 6045 6856
rect 6011 6754 6045 6788
rect 6011 6702 6045 6720
rect 6187 7016 6221 7050
rect 6187 6890 6221 6982
rect 6187 6822 6221 6856
rect 6187 6780 6221 6788
rect 6187 6708 6221 6720
rect 3871 6601 3883 6635
rect 3929 6601 3955 6635
rect 3997 6601 4027 6635
rect 4065 6601 4099 6635
rect 4133 6601 4167 6635
rect 4205 6601 4235 6635
rect 4277 6601 4303 6635
rect 4349 6601 4371 6635
rect 4421 6601 4439 6635
rect 4493 6601 4507 6635
rect 4565 6601 4575 6635
rect 4637 6601 4643 6635
rect 4709 6601 4711 6635
rect 4745 6601 4747 6635
rect 4813 6601 4819 6635
rect 4881 6601 4891 6635
rect 4949 6601 4963 6635
rect 5017 6601 5035 6635
rect 5085 6601 5107 6635
rect 5153 6601 5179 6635
rect 5221 6601 5251 6635
rect 5289 6601 5323 6635
rect 5357 6601 5391 6635
rect 5429 6601 5459 6635
rect 5501 6601 5527 6635
rect 5573 6601 5595 6635
rect 5645 6601 5663 6635
rect 5717 6601 5731 6635
rect 5789 6601 5799 6635
rect 5861 6601 5867 6635
rect 5933 6601 5935 6635
rect 5969 6601 5971 6635
rect 6037 6601 6043 6635
rect 6105 6601 6115 6635
rect 6173 6601 6229 6635
rect 3879 6516 3913 6562
rect 3879 6448 3913 6482
rect 3879 6380 3913 6414
rect 3879 6254 3913 6346
rect 3879 6186 3913 6220
rect 3879 6118 3913 6152
rect 4055 6516 4089 6532
rect 4055 6448 4089 6482
rect 4055 6380 4089 6414
rect 4055 6254 4089 6346
rect 4231 6516 4265 6528
rect 4231 6448 4265 6456
rect 4231 6380 4265 6414
rect 4055 6186 4089 6220
rect 4055 6136 4089 6152
rect 4127 6337 4193 6341
rect 4127 6303 4140 6337
rect 4174 6303 4193 6337
rect 4127 6265 4193 6303
rect 4127 6231 4140 6265
rect 4174 6231 4193 6265
rect 3913 6084 4055 6102
rect 3879 6068 4055 6084
rect 4055 6030 4089 6068
rect 3949 6017 3965 6018
rect 3949 5983 3962 6017
rect 3999 5984 4015 6018
rect 3996 5983 4015 5984
rect 3949 5950 4015 5983
rect 3949 5945 3965 5950
rect 3949 5911 3962 5945
rect 3999 5916 4015 5950
rect 3996 5911 4015 5916
rect 3949 5898 4015 5911
rect 3879 5856 3913 5872
rect 3879 5811 3913 5822
rect 3879 5739 3913 5754
rect 4055 5856 4089 5996
rect 4127 6018 4193 6231
rect 4231 6254 4265 6346
rect 4231 6186 4265 6220
rect 4231 6118 4265 6152
rect 4231 6068 4265 6084
rect 4355 6516 4389 6528
rect 4355 6448 4389 6456
rect 4355 6380 4389 6414
rect 4355 6254 4389 6346
rect 4531 6516 4565 6534
rect 4531 6448 4565 6482
rect 4531 6380 4565 6414
rect 4531 6254 4565 6346
rect 4355 6186 4389 6220
rect 4355 6118 4389 6152
rect 4355 6068 4389 6084
rect 4430 6212 4439 6238
rect 4473 6212 4496 6238
rect 4430 6174 4496 6212
rect 4430 6140 4439 6174
rect 4473 6140 4496 6174
rect 4127 5984 4143 6018
rect 4177 5984 4193 6018
rect 4127 5950 4193 5984
rect 4127 5916 4143 5950
rect 4177 5916 4193 5950
rect 4430 6018 4496 6140
rect 4430 5984 4446 6018
rect 4480 5984 4496 6018
rect 4430 5950 4496 5984
rect 4430 5916 4446 5950
rect 4480 5916 4496 5950
rect 4531 6186 4565 6220
rect 4531 6118 4565 6152
rect 4055 5788 4089 5822
rect 4055 5738 4089 5754
rect 4231 5856 4265 5872
rect 4231 5811 4265 5822
rect 4231 5739 4265 5754
rect 4355 5856 4389 5872
rect 4355 5811 4389 5822
rect 4531 5845 4565 6084
rect 4707 6516 4741 6528
rect 4707 6448 4741 6456
rect 4707 6380 4741 6414
rect 4707 6254 4741 6346
rect 4707 6186 4741 6220
rect 4707 6118 4741 6152
rect 4707 6068 4741 6084
rect 4831 6516 4865 6528
rect 4831 6448 4865 6456
rect 4831 6380 4865 6414
rect 4831 6254 4865 6346
rect 4831 6186 4865 6220
rect 4831 6118 4865 6152
rect 4831 6068 4865 6084
rect 5007 6516 5041 6534
rect 5007 6448 5041 6482
rect 5007 6380 5041 6414
rect 5007 6254 5041 6346
rect 5007 6186 5041 6187
rect 5007 6149 5041 6152
rect 5183 6516 5217 6528
rect 5183 6448 5217 6456
rect 5183 6380 5217 6414
rect 5359 6516 5393 6534
rect 5359 6448 5393 6482
rect 5359 6380 5393 6414
rect 5183 6254 5217 6346
rect 5183 6186 5217 6220
rect 4601 5985 4617 6018
rect 4601 5951 4615 5985
rect 4651 5984 4667 6018
rect 4905 5990 4921 6018
rect 4955 5990 4971 6018
rect 4649 5951 4667 5984
rect 4601 5950 4667 5951
rect 4601 5916 4617 5950
rect 4651 5916 4667 5950
rect 4741 5956 4779 5990
rect 4813 5956 4865 5990
rect 4899 5984 4921 5990
rect 4899 5956 4937 5984
rect 4615 5913 4649 5916
rect 4707 5856 4741 5956
rect 4905 5950 4971 5956
rect 4905 5916 4921 5950
rect 4955 5916 4971 5950
rect 4531 5822 4707 5845
rect 4531 5811 4741 5822
rect 4355 5739 4389 5754
rect 4702 5788 4741 5811
rect 4702 5754 4707 5788
rect 4702 5738 4741 5754
rect 4831 5856 4865 5872
rect 5007 5845 5041 6084
rect 5076 6109 5093 6143
rect 5127 6109 5142 6143
rect 5076 6071 5142 6109
rect 5076 6037 5093 6071
rect 5127 6037 5142 6071
rect 5183 6118 5217 6152
rect 5183 6068 5217 6084
rect 5258 6330 5324 6348
rect 5258 6296 5274 6330
rect 5308 6296 5324 6330
rect 5258 6258 5324 6296
rect 5258 6224 5274 6258
rect 5308 6224 5324 6258
rect 5076 6018 5142 6037
rect 5076 5984 5092 6018
rect 5126 5984 5142 6018
rect 5076 5950 5142 5984
rect 5076 5916 5092 5950
rect 5126 5916 5142 5950
rect 5258 6018 5324 6224
rect 5258 5984 5274 6018
rect 5308 5984 5324 6018
rect 5258 5950 5324 5984
rect 5258 5916 5274 5950
rect 5308 5916 5324 5950
rect 5359 6254 5393 6346
rect 5359 6186 5393 6220
rect 5359 6143 5393 6152
rect 5359 6071 5393 6084
rect 5535 6516 5569 6528
rect 5535 6448 5569 6456
rect 5535 6380 5569 6414
rect 5535 6254 5569 6346
rect 5535 6186 5569 6220
rect 5535 6118 5569 6152
rect 5535 6068 5569 6084
rect 5659 6516 5693 6534
rect 5659 6448 5693 6482
rect 5659 6380 5693 6414
rect 5659 6254 5693 6346
rect 5659 6186 5693 6220
rect 5659 6118 5693 6141
rect 4865 5822 5041 5845
rect 4831 5811 5041 5822
rect 5183 5856 5217 5872
rect 5183 5811 5217 5822
rect 5359 5845 5393 6037
rect 5429 5984 5445 6018
rect 5479 5987 5495 6018
rect 5429 5953 5446 5984
rect 5480 5953 5495 5987
rect 5429 5950 5495 5953
rect 5429 5916 5445 5950
rect 5479 5916 5495 5950
rect 5446 5915 5480 5916
rect 5535 5856 5569 5872
rect 5359 5822 5535 5845
rect 5359 5811 5569 5822
rect 4831 5788 4870 5811
rect 4865 5754 4870 5788
rect 4831 5738 4870 5754
rect 5183 5739 5217 5754
rect 5530 5788 5569 5811
rect 5530 5754 5535 5788
rect 5530 5738 5569 5754
rect 5659 5856 5693 6069
rect 5835 6516 5869 6528
rect 5835 6448 5869 6456
rect 5835 6380 5869 6414
rect 5835 6254 5869 6346
rect 5835 6186 5869 6220
rect 6011 6516 6045 6534
rect 6011 6448 6045 6482
rect 6011 6380 6045 6414
rect 6011 6308 6045 6346
rect 6011 6254 6045 6274
rect 5835 6118 5869 6152
rect 5835 6068 5869 6084
rect 5903 6175 5968 6193
rect 5903 6141 5917 6175
rect 5951 6141 5968 6175
rect 5903 6103 5968 6141
rect 5903 6069 5917 6103
rect 5951 6069 5968 6103
rect 5903 6018 5968 6069
rect 6011 6186 6045 6220
rect 6187 6516 6221 6528
rect 6187 6448 6221 6456
rect 6187 6380 6221 6414
rect 6187 6254 6221 6346
rect 6011 6118 6045 6152
rect 5730 5988 5737 6018
rect 5730 5984 5746 5988
rect 5780 5984 5796 6018
rect 5730 5950 5796 5984
rect 5730 5916 5737 5950
rect 5780 5916 5796 5950
rect 5901 5984 5917 6018
rect 5951 5984 5967 6018
rect 5901 5950 5967 5984
rect 5901 5916 5917 5950
rect 5951 5916 5967 5950
rect 5659 5788 5693 5822
rect 5659 5738 5693 5754
rect 5835 5856 5869 5872
rect 5835 5811 5869 5822
rect 5835 5739 5869 5754
rect 6011 5856 6045 6084
rect 6089 6175 6152 6193
rect 6089 6141 6111 6175
rect 6145 6141 6152 6175
rect 6089 6103 6152 6141
rect 6089 6069 6111 6103
rect 6145 6069 6152 6103
rect 6089 6018 6152 6069
rect 6187 6186 6221 6220
rect 6187 6118 6221 6152
rect 6187 6068 6221 6084
rect 6088 5984 6104 6018
rect 6138 5984 6154 6018
rect 6088 5950 6154 5984
rect 6088 5916 6104 5950
rect 6138 5916 6154 5950
rect 6011 5788 6045 5822
rect 6011 5738 6045 5754
rect 6187 5856 6221 5872
rect 6187 5811 6221 5822
rect 6187 5739 6221 5754
rect 3868 5620 3880 5654
rect 3926 5620 3952 5654
rect 3994 5620 4024 5654
rect 4062 5620 4096 5654
rect 4130 5620 4164 5654
rect 4202 5620 4232 5654
rect 4274 5620 4300 5654
rect 4346 5620 4368 5654
rect 4418 5620 4436 5654
rect 4490 5620 4504 5654
rect 4562 5620 4572 5654
rect 4634 5620 4640 5654
rect 4706 5620 4708 5654
rect 4742 5620 4744 5654
rect 4810 5620 4816 5654
rect 4878 5620 4888 5654
rect 4946 5620 4960 5654
rect 5014 5620 5032 5654
rect 5082 5620 5104 5654
rect 5150 5620 5176 5654
rect 5218 5620 5248 5654
rect 5286 5620 5320 5654
rect 5354 5620 5388 5654
rect 5426 5620 5456 5654
rect 5498 5620 5524 5654
rect 5570 5620 5592 5654
rect 5642 5620 5660 5654
rect 5714 5620 5728 5654
rect 5786 5620 5796 5654
rect 5858 5620 5864 5654
rect 5930 5620 5932 5654
rect 5966 5620 5968 5654
rect 6034 5620 6040 5654
rect 6102 5620 6112 5654
rect 6170 5620 6184 5654
rect 6218 5620 6254 5654
rect 5324 5581 6254 5620
rect 4019 5531 4035 5565
rect 4069 5531 4112 5565
rect 4146 5531 4189 5565
rect 4223 5531 4265 5565
rect 4299 5531 4315 5565
rect 4363 5531 4379 5565
rect 4413 5531 4447 5565
rect 4481 5531 4907 5565
rect 4941 5531 4975 5565
rect 5009 5531 5025 5565
rect 5324 5547 5336 5581
rect 5382 5547 5408 5581
rect 5450 5547 5480 5581
rect 5518 5547 5552 5581
rect 5586 5547 5620 5581
rect 5658 5547 5688 5581
rect 5730 5547 5756 5581
rect 5802 5547 5824 5581
rect 5874 5547 5892 5581
rect 5946 5547 5960 5581
rect 6018 5547 6028 5581
rect 6090 5547 6096 5581
rect 6162 5547 6164 5581
rect 6198 5547 6200 5581
rect 6234 5547 6254 5581
rect 3974 5477 4008 5493
rect 3974 5409 4008 5443
rect 3974 5172 4008 5375
rect 4150 5477 4184 5493
rect 4150 5409 4184 5435
rect 4150 5359 4184 5363
rect 4218 5317 4292 5531
rect 4326 5477 4360 5493
rect 4326 5409 4360 5443
rect 4326 5359 4360 5375
rect 4502 5477 4536 5493
rect 4502 5409 4536 5443
rect 4233 5283 4271 5317
rect 4008 5138 4046 5172
rect 3974 5075 4008 5138
rect 3974 5007 4008 5041
rect 3974 4939 4008 4973
rect 3974 4807 4008 4905
rect 3974 4739 4008 4773
rect 3974 4671 4008 4705
rect 3974 4621 4008 4637
rect 4150 5075 4184 5091
rect 4150 5007 4184 5041
rect 4150 4939 4184 4973
rect 4150 4807 4184 4905
rect 4150 4739 4184 4773
rect 4150 4671 4184 4703
rect 4150 4621 4184 4631
rect 4218 4571 4292 5283
rect 4413 5249 4447 5263
rect 4396 5247 4434 5249
rect 4396 5215 4413 5247
rect 4413 5179 4447 5213
rect 4413 5129 4447 5145
rect 4326 5075 4360 5091
rect 4326 5007 4360 5041
rect 4326 4939 4360 4973
rect 4326 4807 4360 4905
rect 4502 5075 4536 5375
rect 4678 5477 4712 5493
rect 4678 5409 4712 5443
rect 4678 5359 4712 5375
rect 4502 5007 4536 5041
rect 4502 4939 4536 4973
rect 4502 4836 4536 4905
rect 4463 4802 4501 4836
rect 4535 4807 4536 4836
rect 4326 4739 4360 4773
rect 4326 4671 4360 4705
rect 4326 4621 4360 4637
rect 4502 4739 4536 4773
rect 4502 4671 4536 4705
rect 4502 4621 4536 4637
rect 4570 5172 4644 5174
rect 4604 5138 4642 5172
rect 4570 4571 4644 5138
rect 4678 5075 4712 5091
rect 4678 5007 4712 5041
rect 4678 4939 4712 4973
rect 4678 4807 4712 4905
rect 4678 4739 4712 4773
rect 4678 4671 4712 4705
rect 4678 4621 4712 4637
rect 4746 4977 4820 5531
rect 5324 5507 6254 5547
rect 4854 5477 4888 5493
rect 4854 5409 4888 5435
rect 4854 5359 4888 5363
rect 5030 5477 5064 5493
rect 5324 5473 5336 5507
rect 5382 5473 5408 5507
rect 5450 5473 5480 5507
rect 5518 5473 5552 5507
rect 5586 5473 5620 5507
rect 5658 5473 5688 5507
rect 5730 5473 5756 5507
rect 5802 5473 5824 5507
rect 5874 5473 5892 5507
rect 5946 5473 5960 5507
rect 6018 5473 6028 5507
rect 6090 5473 6096 5507
rect 6162 5473 6164 5507
rect 6198 5473 6200 5507
rect 6234 5473 6254 5507
rect 5030 5409 5064 5443
rect 5030 5249 5064 5375
rect 4992 5215 5030 5249
rect 5348 5356 5382 5371
rect 5348 5288 5382 5299
rect 5348 5238 5382 5254
rect 5524 5356 5558 5372
rect 5524 5288 5558 5322
rect 4746 4943 4766 4977
rect 4800 4943 4820 4977
rect 4746 4905 4820 4943
rect 4746 4871 4766 4905
rect 4800 4871 4820 4905
rect 4746 4571 4820 4871
rect 4854 5075 4888 5091
rect 4854 5007 4888 5041
rect 4854 4939 4888 4973
rect 4854 4807 4888 4905
rect 4854 4739 4888 4773
rect 4854 4671 4888 4703
rect 4854 4621 4888 4631
rect 5030 5075 5064 5215
rect 5421 5160 5437 5194
rect 5471 5160 5487 5194
rect 5421 5126 5487 5160
rect 5421 5092 5437 5126
rect 5471 5092 5487 5126
rect 5421 5045 5487 5092
rect 5030 5007 5064 5041
rect 5030 4939 5064 4973
rect 5030 4807 5064 4905
rect 5030 4739 5064 4773
rect 5030 4671 5064 4705
rect 5030 4621 5064 4637
rect 5348 5026 5382 5042
rect 5348 4958 5382 4992
rect 5421 5011 5435 5045
rect 5469 5011 5487 5045
rect 5421 4973 5487 5011
rect 5421 4939 5435 4973
rect 5469 4939 5487 4973
rect 5524 5156 5558 5254
rect 5648 5356 5682 5371
rect 5648 5288 5682 5299
rect 5648 5238 5682 5254
rect 5824 5356 5858 5372
rect 5824 5288 5858 5322
rect 5524 5084 5558 5122
rect 5715 5160 5731 5194
rect 5765 5160 5781 5194
rect 5715 5126 5781 5160
rect 5715 5092 5731 5126
rect 5765 5092 5781 5126
rect 5524 5026 5558 5050
rect 5524 4958 5558 4992
rect 5348 4890 5382 4924
rect 5348 4764 5382 4856
rect 5348 4696 5382 4730
rect 5348 4654 5382 4662
rect 5348 4582 5382 4594
rect 4019 4537 4035 4571
rect 4069 4537 4112 4571
rect 4146 4537 4189 4571
rect 4223 4537 4265 4571
rect 4299 4537 4315 4571
rect 4539 4537 4555 4571
rect 4589 4537 4623 4571
rect 4657 4537 4673 4571
rect 4723 4537 4739 4571
rect 4773 4537 4816 4571
rect 4850 4537 4893 4571
rect 4927 4537 4969 4571
rect 5003 4537 5019 4571
rect 5524 4890 5558 4924
rect 5524 4764 5558 4856
rect 5524 4696 5558 4730
rect 5524 4628 5558 4662
rect 5524 4576 5558 4594
rect 5648 5026 5682 5042
rect 5648 4958 5682 4992
rect 5648 4890 5682 4924
rect 5716 5041 5781 5092
rect 5716 5007 5725 5041
rect 5759 5007 5781 5041
rect 5716 4969 5781 5007
rect 5716 4935 5725 4969
rect 5759 4935 5781 4969
rect 5716 4917 5781 4935
rect 5824 5026 5858 5254
rect 6000 5356 6034 5371
rect 6000 5288 6034 5299
rect 6000 5238 6034 5254
rect 6176 5356 6210 5372
rect 6176 5288 6210 5322
rect 5824 4958 5858 4992
rect 5648 4764 5682 4856
rect 5824 4890 5858 4924
rect 5902 5160 5918 5194
rect 5952 5160 5968 5194
rect 5902 5126 5968 5160
rect 5902 5092 5918 5126
rect 5952 5092 5968 5126
rect 6073 5170 6088 5194
rect 6073 5160 6089 5170
rect 6123 5160 6139 5194
rect 6073 5132 6139 5160
rect 6073 5098 6088 5132
rect 6122 5126 6139 5132
rect 6073 5092 6089 5098
rect 6123 5092 6139 5126
rect 5902 5041 5966 5092
rect 5902 5007 5919 5041
rect 5953 5007 5966 5041
rect 5902 4969 5966 5007
rect 5902 4935 5919 4969
rect 5953 4935 5966 4969
rect 5902 4917 5966 4935
rect 6000 5026 6034 5042
rect 6000 4958 6034 4992
rect 5824 4834 5858 4856
rect 5648 4696 5682 4730
rect 5857 4800 5858 4834
rect 5823 4764 5858 4800
rect 5823 4762 5824 4764
rect 5857 4728 5858 4730
rect 5648 4654 5682 4662
rect 5648 4582 5682 4594
rect 5824 4696 5858 4728
rect 5824 4628 5858 4662
rect 5824 4576 5858 4594
rect 6000 4890 6034 4924
rect 6000 4764 6034 4856
rect 6000 4696 6034 4730
rect 6000 4654 6034 4662
rect 6000 4582 6034 4594
rect 6176 5041 6210 5254
rect 6176 5026 6177 5041
rect 6210 4992 6211 5007
rect 6176 4969 6211 4992
rect 6176 4958 6177 4969
rect 6176 4890 6210 4924
rect 6176 4764 6210 4856
rect 6176 4696 6210 4730
rect 6176 4628 6210 4662
rect 6176 4576 6210 4594
rect 5194 4470 5230 4501
rect 3996 4436 4035 4470
rect 4089 4436 4103 4470
rect 4161 4436 4171 4470
rect 4233 4436 4239 4470
rect 4305 4436 4307 4470
rect 4341 4436 4343 4470
rect 4409 4436 4415 4470
rect 4477 4436 4487 4470
rect 4545 4436 4559 4470
rect 4613 4436 4631 4470
rect 4681 4436 4703 4470
rect 4749 4436 4775 4470
rect 4817 4436 4847 4470
rect 4885 4436 4919 4470
rect 4953 4436 4987 4470
rect 5025 4436 5055 4470
rect 5097 4436 5123 4470
rect 5169 4467 5230 4470
rect 5264 4467 5298 4501
rect 5336 4467 5366 4501
rect 5408 4467 5434 4501
rect 5480 4467 5502 4501
rect 5552 4467 5570 4501
rect 5624 4467 5638 4501
rect 5696 4467 5706 4501
rect 5768 4467 5774 4501
rect 5840 4467 5842 4501
rect 5876 4467 5878 4501
rect 5944 4467 5950 4501
rect 6012 4467 6022 4501
rect 6080 4467 6094 4501
rect 6148 4467 6218 4501
rect 5169 4436 5228 4467
rect 5323 4374 5357 4420
rect 3986 4332 4002 4366
rect 4036 4332 4079 4366
rect 4113 4332 4156 4366
rect 4190 4332 4232 4366
rect 4266 4332 4282 4366
rect 4506 4332 4522 4366
rect 4556 4332 4590 4366
rect 4624 4332 4640 4366
rect 4690 4332 4706 4366
rect 4740 4332 4783 4366
rect 4817 4332 4860 4366
rect 4894 4332 4936 4366
rect 4970 4332 4986 4366
rect 3941 4266 3975 4282
rect 3941 4198 3975 4232
rect 3941 4130 3975 4164
rect 3941 3998 3975 4096
rect 3941 3930 3975 3964
rect 3941 3862 3975 3896
rect 3941 3765 3975 3828
rect 4117 4272 4151 4282
rect 4117 4200 4151 4232
rect 4117 4130 4151 4164
rect 4117 3998 4151 4096
rect 4117 3930 4151 3964
rect 4117 3862 4151 3896
rect 4117 3812 4151 3828
rect 4185 3956 4259 4332
rect 4185 3922 4199 3956
rect 4233 3922 4259 3956
rect 4185 3884 4259 3922
rect 4185 3850 4199 3884
rect 4233 3850 4259 3884
rect 3975 3731 4013 3765
rect 3941 3528 3975 3731
rect 3941 3460 3975 3494
rect 3941 3410 3975 3426
rect 4117 3540 4151 3544
rect 4117 3468 4151 3494
rect 4117 3410 4151 3426
rect 4185 3372 4259 3850
rect 4293 4266 4327 4282
rect 4293 4198 4327 4232
rect 4293 4130 4327 4164
rect 4293 3998 4327 4096
rect 4469 4266 4503 4282
rect 4469 4198 4503 4232
rect 4469 4130 4503 4164
rect 4469 3998 4503 4096
rect 4293 3930 4327 3964
rect 4429 3935 4467 3969
rect 4501 3935 4503 3964
rect 4293 3862 4327 3896
rect 4293 3812 4327 3828
rect 4469 3930 4503 3935
rect 4469 3862 4503 3896
rect 4380 3758 4414 3774
rect 4380 3690 4414 3724
rect 4363 3656 4380 3688
rect 4363 3654 4401 3656
rect 4380 3640 4414 3654
rect 4293 3528 4327 3544
rect 4293 3460 4327 3494
rect 4293 3410 4327 3426
rect 4469 3528 4503 3828
rect 4537 3765 4611 4332
rect 4645 4266 4679 4282
rect 4645 4198 4679 4232
rect 4645 4130 4679 4164
rect 4645 3998 4679 4096
rect 4645 3930 4679 3964
rect 4645 3862 4679 3896
rect 4645 3812 4679 3828
rect 4713 3869 4787 4332
rect 5323 4306 5357 4340
rect 4713 3835 4736 3869
rect 4770 3835 4787 3869
rect 4713 3797 4787 3835
rect 4821 4272 4855 4282
rect 4821 4200 4855 4232
rect 4821 4130 4855 4164
rect 4821 3998 4855 4096
rect 4821 3930 4855 3964
rect 4821 3862 4855 3896
rect 4821 3812 4855 3828
rect 4997 4266 5031 4282
rect 4997 4198 5031 4232
rect 4997 4130 5031 4164
rect 4997 3998 5031 4096
rect 4997 3930 5031 3964
rect 5323 4246 5357 4272
rect 5323 4174 5357 4204
rect 5323 4112 5357 4140
rect 5323 4044 5357 4078
rect 5323 3976 5357 4010
rect 5499 4374 5533 4390
rect 5499 4306 5533 4340
rect 5499 4238 5533 4272
rect 5499 4112 5533 4204
rect 5499 4044 5533 4078
rect 5499 3994 5533 4010
rect 5675 4374 5709 4386
rect 5675 4306 5709 4314
rect 5675 4238 5709 4272
rect 5675 4112 5709 4204
rect 5675 4044 5709 4078
rect 5851 4374 5885 4392
rect 5851 4306 5885 4340
rect 5851 4238 5885 4272
rect 5851 4112 5885 4204
rect 5675 3976 5709 4010
rect 5357 3942 5533 3960
rect 5323 3926 5533 3942
rect 5675 3926 5709 3942
rect 5744 4033 5808 4049
rect 5744 3999 5752 4033
rect 5786 3999 5808 4033
rect 5744 3961 5808 3999
rect 5744 3927 5752 3961
rect 5786 3927 5808 3961
rect 4997 3862 5031 3896
rect 4571 3731 4609 3765
rect 4537 3709 4643 3731
rect 4713 3763 4736 3797
rect 4770 3763 4787 3797
rect 4537 3675 4553 3709
rect 4587 3675 4621 3709
rect 4655 3675 4671 3709
rect 4469 3460 4503 3494
rect 4469 3410 4503 3426
rect 4645 3528 4679 3544
rect 4645 3460 4679 3494
rect 4645 3410 4679 3426
rect 4713 3372 4787 3763
rect 4997 3688 5031 3828
rect 5393 3842 5409 3876
rect 5443 3842 5459 3876
rect 5393 3808 5459 3842
rect 5393 3774 5409 3808
rect 5443 3774 5459 3808
rect 4959 3654 4997 3688
rect 4821 3540 4855 3544
rect 4821 3468 4855 3494
rect 4821 3410 4855 3426
rect 4997 3528 5031 3654
rect 5323 3714 5357 3730
rect 5323 3669 5357 3680
rect 5323 3597 5357 3612
rect 5499 3714 5533 3926
rect 5744 3876 5808 3927
rect 5851 4044 5885 4078
rect 6027 4374 6061 4386
rect 6027 4306 6061 4314
rect 6027 4238 6061 4272
rect 6203 4374 6237 4392
rect 6203 4306 6237 4340
rect 6027 4112 6061 4204
rect 5851 3976 5885 4010
rect 5851 3885 5885 3942
rect 5571 3842 5587 3876
rect 5622 3842 5637 3876
rect 5571 3808 5637 3842
rect 5571 3774 5587 3808
rect 5621 3804 5637 3808
rect 5622 3774 5637 3804
rect 5742 3842 5758 3876
rect 5792 3842 5808 3876
rect 5742 3808 5808 3842
rect 5742 3774 5758 3808
rect 5792 3774 5808 3808
rect 5884 3851 5885 3885
rect 5850 3813 5885 3851
rect 5884 3779 5885 3813
rect 5499 3646 5533 3680
rect 5499 3596 5533 3612
rect 5675 3714 5709 3730
rect 5675 3669 5709 3680
rect 5675 3597 5709 3612
rect 5851 3714 5885 3779
rect 5929 4031 5992 4049
rect 5929 3997 5946 4031
rect 5980 3997 5992 4031
rect 5929 3959 5992 3997
rect 5929 3925 5946 3959
rect 5980 3925 5992 3959
rect 6027 4044 6061 4078
rect 6027 3976 6061 4010
rect 6027 3926 6061 3942
rect 6100 4212 6116 4246
rect 6150 4212 6166 4246
rect 6100 4174 6166 4212
rect 6100 4140 6116 4174
rect 6150 4140 6166 4174
rect 5929 3876 5992 3925
rect 6100 3876 6166 4140
rect 5929 3842 5945 3876
rect 5979 3842 5995 3876
rect 5929 3808 5995 3842
rect 5929 3774 5945 3808
rect 5979 3774 5995 3808
rect 6100 3842 6116 3876
rect 6150 3842 6166 3876
rect 6100 3808 6166 3842
rect 6100 3774 6116 3808
rect 6150 3774 6166 3808
rect 6203 4238 6237 4272
rect 6203 4112 6237 4204
rect 6203 4044 6237 4078
rect 6203 3997 6204 4010
rect 6203 3976 6238 3997
rect 6237 3959 6238 3976
rect 6203 3925 6204 3942
rect 5851 3646 5885 3680
rect 5851 3596 5885 3612
rect 6027 3714 6061 3730
rect 6027 3669 6061 3680
rect 6027 3597 6061 3612
rect 6203 3714 6237 3925
rect 6203 3646 6237 3680
rect 6203 3596 6237 3612
rect 4997 3460 5031 3494
rect 4997 3410 5031 3426
rect 5114 3478 5126 3512
rect 5172 3478 5198 3512
rect 5240 3478 5270 3512
rect 5308 3478 5342 3512
rect 5376 3478 5410 3512
rect 5448 3478 5478 3512
rect 5520 3478 5546 3512
rect 5592 3478 5614 3512
rect 5664 3478 5682 3512
rect 5736 3478 5750 3512
rect 5808 3478 5818 3512
rect 5880 3478 5886 3512
rect 5952 3478 5954 3512
rect 5988 3478 5990 3512
rect 6056 3478 6062 3512
rect 6124 3478 6134 3512
rect 6192 3478 6206 3512
rect 6240 3478 6265 3512
rect 5114 3444 5148 3478
rect 5114 3384 5148 3410
rect 3986 3338 4002 3372
rect 4036 3338 4079 3372
rect 4113 3338 4156 3372
rect 4190 3338 4232 3372
rect 4266 3338 4282 3372
rect 4330 3338 4346 3372
rect 4380 3338 4414 3372
rect 4448 3338 4874 3372
rect 4908 3338 4942 3372
rect 4976 3338 4992 3372
rect -9272 2834 -9238 2880
rect -9272 2766 -9238 2800
rect -9272 2698 -9238 2732
rect -9272 2572 -9238 2664
rect -9272 2504 -9238 2538
rect -9272 2436 -9238 2470
rect -9096 2834 -9062 2850
rect -9096 2766 -9062 2800
rect -9096 2698 -9062 2732
rect -9096 2572 -9062 2664
rect -9096 2504 -9062 2538
rect -8920 2834 -8886 2846
rect -8920 2766 -8886 2774
rect -8920 2698 -8886 2732
rect -8920 2572 -8886 2664
rect -8920 2504 -8886 2538
rect -9096 2454 -9062 2470
rect -9024 2453 -9006 2487
rect -8972 2453 -8958 2487
rect -9238 2402 -9062 2420
rect -9272 2386 -9062 2402
rect -9202 2336 -9180 2343
rect -9202 2302 -9186 2336
rect -9146 2309 -9136 2343
rect -9152 2302 -9136 2309
rect -9202 2271 -9136 2302
rect -9202 2268 -9180 2271
rect -9202 2234 -9186 2268
rect -9146 2237 -9136 2271
rect -9152 2234 -9136 2237
rect -9096 2336 -9062 2386
rect -9096 2264 -9062 2302
rect -9024 2415 -8958 2453
rect -9024 2381 -9006 2415
rect -8972 2381 -8958 2415
rect -8744 2834 -8710 2852
rect -8744 2766 -8710 2800
rect -8744 2698 -8710 2732
rect -8744 2572 -8710 2664
rect -8744 2533 -8710 2538
rect -8920 2436 -8886 2470
rect -8920 2386 -8886 2402
rect -8845 2453 -8827 2487
rect -8793 2453 -8779 2487
rect -8845 2415 -8779 2453
rect -9024 2336 -8958 2381
rect -9024 2302 -9008 2336
rect -8974 2302 -8958 2336
rect -9024 2268 -8958 2302
rect -9024 2234 -9008 2268
rect -8974 2234 -8958 2268
rect -8845 2381 -8827 2415
rect -8793 2381 -8779 2415
rect -8845 2336 -8779 2381
rect -8845 2302 -8829 2336
rect -8795 2302 -8779 2336
rect -8845 2268 -8779 2302
rect -8845 2234 -8829 2268
rect -8795 2234 -8779 2268
rect -8744 2461 -8710 2470
rect -9272 2174 -9238 2190
rect -9272 2129 -9238 2140
rect -9272 2057 -9238 2072
rect -9096 2174 -9062 2230
rect -9096 2106 -9062 2140
rect -9096 2056 -9062 2072
rect -8920 2174 -8886 2190
rect -8920 2129 -8886 2140
rect -8744 2163 -8710 2402
rect -8568 2834 -8534 2846
rect -8568 2766 -8534 2774
rect -8568 2698 -8534 2732
rect -8568 2572 -8534 2664
rect -8568 2504 -8534 2538
rect -8568 2436 -8534 2470
rect -8568 2386 -8534 2402
rect -8674 2302 -8658 2336
rect -8615 2302 -8608 2336
rect -8674 2268 -8608 2302
rect -8674 2234 -8658 2268
rect -8624 2264 -8608 2268
rect -8615 2234 -8608 2264
rect -8568 2174 -8534 2190
rect -8744 2140 -8568 2163
rect -8744 2129 -8534 2140
rect -8920 2057 -8886 2072
rect -8573 2106 -8534 2129
rect -8573 2072 -8568 2106
rect -8573 2056 -8534 2072
<< viali >>
rect 3883 7582 3895 7616
rect 3895 7582 3917 7616
rect 3955 7582 3963 7616
rect 3963 7582 3989 7616
rect 4027 7582 4031 7616
rect 4031 7582 4061 7616
rect 4099 7582 4133 7616
rect 4171 7582 4201 7616
rect 4201 7582 4205 7616
rect 4243 7582 4269 7616
rect 4269 7582 4277 7616
rect 4315 7582 4337 7616
rect 4337 7582 4349 7616
rect 4387 7582 4405 7616
rect 4405 7582 4421 7616
rect 4459 7582 4473 7616
rect 4473 7582 4493 7616
rect 4531 7582 4541 7616
rect 4541 7582 4565 7616
rect 4603 7582 4609 7616
rect 4609 7582 4637 7616
rect 4675 7582 4677 7616
rect 4677 7582 4709 7616
rect 4747 7582 4779 7616
rect 4779 7582 4781 7616
rect 4819 7582 4847 7616
rect 4847 7582 4853 7616
rect 4891 7582 4915 7616
rect 4915 7582 4925 7616
rect 4963 7582 4983 7616
rect 4983 7582 4997 7616
rect 5035 7582 5051 7616
rect 5051 7582 5069 7616
rect 5107 7582 5119 7616
rect 5119 7582 5141 7616
rect 5179 7582 5187 7616
rect 5187 7582 5213 7616
rect 5251 7582 5255 7616
rect 5255 7582 5285 7616
rect 5323 7582 5357 7616
rect 5395 7582 5425 7616
rect 5425 7582 5429 7616
rect 5467 7582 5493 7616
rect 5493 7582 5501 7616
rect 5539 7582 5561 7616
rect 5561 7582 5573 7616
rect 5611 7582 5629 7616
rect 5629 7582 5645 7616
rect 5683 7582 5697 7616
rect 5697 7582 5717 7616
rect 5755 7582 5765 7616
rect 5765 7582 5789 7616
rect 5827 7582 5833 7616
rect 5833 7582 5861 7616
rect 5899 7582 5901 7616
rect 5901 7582 5933 7616
rect 5971 7582 6003 7616
rect 6003 7582 6005 7616
rect 6043 7582 6071 7616
rect 6071 7582 6077 7616
rect 6115 7582 6139 7616
rect 6139 7582 6149 7616
rect 6187 7582 6221 7616
rect 4231 7497 4265 7531
rect 4231 7448 4265 7459
rect 4231 7425 4265 7448
rect 3971 7286 4003 7302
rect 4003 7286 4005 7302
rect 3971 7268 4005 7286
rect 3971 7218 4003 7230
rect 4003 7218 4005 7230
rect 3971 7196 4005 7218
rect 3879 6754 3913 6780
rect 3879 6746 3913 6754
rect 3879 6674 3913 6708
rect 4707 7497 4741 7531
rect 4707 7448 4741 7459
rect 4707 7425 4741 7448
rect 4055 7050 4089 7054
rect 4055 7020 4089 7050
rect 4055 6948 4089 6982
rect 4443 7286 4445 7305
rect 4445 7286 4477 7305
rect 4443 7271 4477 7286
rect 4443 7218 4445 7233
rect 4445 7218 4477 7233
rect 4443 7199 4477 7218
rect 4144 6905 4178 6939
rect 4144 6833 4178 6867
rect 4231 6754 4265 6780
rect 4231 6746 4265 6754
rect 4231 6674 4265 6708
rect 4612 7286 4616 7305
rect 4616 7286 4646 7305
rect 4612 7271 4646 7286
rect 4612 7218 4616 7233
rect 4616 7218 4646 7233
rect 4795 7286 4798 7309
rect 4798 7286 4829 7309
rect 4795 7275 4829 7286
rect 4795 7218 4798 7237
rect 4798 7218 4829 7237
rect 4612 7199 4646 7218
rect 4795 7203 4829 7218
rect 4530 7152 4564 7157
rect 4530 7123 4531 7152
rect 4531 7123 4564 7152
rect 4530 7084 4564 7085
rect 4530 7051 4531 7084
rect 4531 7051 4564 7084
rect 4355 6754 4389 6780
rect 4355 6746 4389 6754
rect 4355 6674 4389 6708
rect 4707 6754 4741 6780
rect 4707 6746 4741 6754
rect 4707 6674 4741 6708
rect 5535 7497 5569 7531
rect 5535 7448 5569 7459
rect 5535 7425 5569 7448
rect 4968 7286 4969 7309
rect 4969 7286 5002 7309
rect 4968 7275 5002 7286
rect 4968 7218 4969 7237
rect 4969 7218 5002 7237
rect 4968 7203 5002 7218
rect 4883 7016 4917 7025
rect 4883 6991 4917 7016
rect 4883 6919 4917 6953
rect 5059 6754 5093 6780
rect 5059 6746 5093 6754
rect 5059 6674 5093 6708
rect 5267 6991 5301 7025
rect 5267 6919 5301 6953
rect 5445 7286 5478 7309
rect 5478 7286 5479 7309
rect 5445 7275 5479 7286
rect 5445 7218 5478 7237
rect 5478 7218 5479 7237
rect 5445 7203 5479 7218
rect 5359 7016 5393 7027
rect 5359 6993 5393 7016
rect 5359 6921 5393 6955
rect 5183 6754 5217 6780
rect 5183 6746 5217 6754
rect 5183 6674 5217 6708
rect 5535 6754 5569 6780
rect 5535 6746 5569 6754
rect 5535 6674 5569 6708
rect 5835 7497 5869 7531
rect 5835 7448 5869 7459
rect 5835 7425 5869 7448
rect 5659 7152 5693 7167
rect 5659 7133 5693 7152
rect 5659 7084 5693 7095
rect 5659 7061 5693 7084
rect 5743 7000 5777 7034
rect 5743 6928 5777 6962
rect 5917 7133 5951 7167
rect 5917 7061 5951 7095
rect 6187 7497 6221 7531
rect 6187 7448 6221 7459
rect 6187 7425 6221 7448
rect 5835 6754 5869 6780
rect 5835 6746 5869 6754
rect 5835 6674 5869 6708
rect 6111 7133 6145 7167
rect 6111 7061 6145 7095
rect 6011 6948 6045 6982
rect 6011 6890 6045 6910
rect 6011 6876 6045 6890
rect 6187 6754 6221 6780
rect 6187 6746 6221 6754
rect 6187 6674 6221 6708
rect 3883 6601 3895 6635
rect 3895 6601 3917 6635
rect 3955 6601 3963 6635
rect 3963 6601 3989 6635
rect 4027 6601 4031 6635
rect 4031 6601 4061 6635
rect 4099 6601 4133 6635
rect 4171 6601 4201 6635
rect 4201 6601 4205 6635
rect 4243 6601 4269 6635
rect 4269 6601 4277 6635
rect 4315 6601 4337 6635
rect 4337 6601 4349 6635
rect 4387 6601 4405 6635
rect 4405 6601 4421 6635
rect 4459 6601 4473 6635
rect 4473 6601 4493 6635
rect 4531 6601 4541 6635
rect 4541 6601 4565 6635
rect 4603 6601 4609 6635
rect 4609 6601 4637 6635
rect 4675 6601 4677 6635
rect 4677 6601 4709 6635
rect 4747 6601 4779 6635
rect 4779 6601 4781 6635
rect 4819 6601 4847 6635
rect 4847 6601 4853 6635
rect 4891 6601 4915 6635
rect 4915 6601 4925 6635
rect 4963 6601 4983 6635
rect 4983 6601 4997 6635
rect 5035 6601 5051 6635
rect 5051 6601 5069 6635
rect 5107 6601 5119 6635
rect 5119 6601 5141 6635
rect 5179 6601 5187 6635
rect 5187 6601 5213 6635
rect 5251 6601 5255 6635
rect 5255 6601 5285 6635
rect 5323 6601 5357 6635
rect 5395 6601 5425 6635
rect 5425 6601 5429 6635
rect 5467 6601 5493 6635
rect 5493 6601 5501 6635
rect 5539 6601 5561 6635
rect 5561 6601 5573 6635
rect 5611 6601 5629 6635
rect 5629 6601 5645 6635
rect 5683 6601 5697 6635
rect 5697 6601 5717 6635
rect 5755 6601 5765 6635
rect 5765 6601 5789 6635
rect 5827 6601 5833 6635
rect 5833 6601 5861 6635
rect 5899 6601 5901 6635
rect 5901 6601 5933 6635
rect 5971 6601 6003 6635
rect 6003 6601 6005 6635
rect 6043 6601 6071 6635
rect 6071 6601 6077 6635
rect 6115 6601 6139 6635
rect 6139 6601 6149 6635
rect 4231 6528 4265 6562
rect 4231 6482 4265 6490
rect 4231 6456 4265 6482
rect 4140 6303 4174 6337
rect 4140 6231 4174 6265
rect 4055 6068 4089 6102
rect 3962 5984 3965 6017
rect 3965 5984 3996 6017
rect 3962 5983 3996 5984
rect 3962 5916 3965 5945
rect 3965 5916 3996 5945
rect 3962 5911 3996 5916
rect 4055 5996 4089 6030
rect 3879 5788 3913 5811
rect 3879 5777 3913 5788
rect 3879 5705 3913 5739
rect 4355 6528 4389 6562
rect 4355 6482 4389 6490
rect 4355 6456 4389 6482
rect 4439 6212 4473 6246
rect 4439 6140 4473 6174
rect 4231 5788 4265 5811
rect 4231 5777 4265 5788
rect 4231 5705 4265 5739
rect 4707 6528 4741 6562
rect 4707 6482 4741 6490
rect 4707 6456 4741 6482
rect 4831 6528 4865 6562
rect 4831 6482 4865 6490
rect 4831 6456 4865 6482
rect 5007 6220 5041 6221
rect 5007 6187 5041 6220
rect 5007 6118 5041 6149
rect 5183 6528 5217 6562
rect 5183 6482 5217 6490
rect 5183 6456 5217 6482
rect 5007 6115 5041 6118
rect 4615 5984 4617 5985
rect 4617 5984 4649 5985
rect 4615 5951 4649 5984
rect 4707 5956 4741 5990
rect 4779 5956 4813 5990
rect 4865 5956 4899 5990
rect 4937 5984 4955 5990
rect 4955 5984 4971 5990
rect 4937 5956 4971 5984
rect 4615 5879 4649 5913
rect 4355 5788 4389 5811
rect 4355 5777 4389 5788
rect 4355 5705 4389 5739
rect 5093 6109 5127 6143
rect 5093 6037 5127 6071
rect 5274 6296 5308 6330
rect 5274 6224 5308 6258
rect 5359 6118 5393 6143
rect 5359 6109 5393 6118
rect 5359 6037 5393 6071
rect 5535 6528 5569 6562
rect 5535 6482 5569 6490
rect 5535 6456 5569 6482
rect 5659 6152 5693 6175
rect 5659 6141 5693 6152
rect 5659 6084 5693 6103
rect 5659 6069 5693 6084
rect 5446 5984 5479 5987
rect 5479 5984 5480 5987
rect 5446 5953 5480 5984
rect 5446 5881 5480 5915
rect 5183 5788 5217 5811
rect 5183 5777 5217 5788
rect 5183 5705 5217 5739
rect 5835 6528 5869 6562
rect 5835 6482 5869 6490
rect 5835 6456 5869 6482
rect 6011 6346 6045 6380
rect 6011 6274 6045 6308
rect 5917 6141 5951 6175
rect 5917 6069 5951 6103
rect 5737 6018 5771 6022
rect 6187 6528 6221 6562
rect 6187 6482 6221 6490
rect 6187 6456 6221 6482
rect 5737 5988 5746 6018
rect 5746 5988 5771 6018
rect 5737 5916 5746 5950
rect 5746 5916 5771 5950
rect 5835 5788 5869 5811
rect 5835 5777 5869 5788
rect 5835 5705 5869 5739
rect 6111 6141 6145 6175
rect 6111 6069 6145 6103
rect 6187 5788 6221 5811
rect 6187 5777 6221 5788
rect 6187 5705 6221 5739
rect 3880 5620 3892 5654
rect 3892 5620 3914 5654
rect 3952 5620 3960 5654
rect 3960 5620 3986 5654
rect 4024 5620 4028 5654
rect 4028 5620 4058 5654
rect 4096 5620 4130 5654
rect 4168 5620 4198 5654
rect 4198 5620 4202 5654
rect 4240 5620 4266 5654
rect 4266 5620 4274 5654
rect 4312 5620 4334 5654
rect 4334 5620 4346 5654
rect 4384 5620 4402 5654
rect 4402 5620 4418 5654
rect 4456 5620 4470 5654
rect 4470 5620 4490 5654
rect 4528 5620 4538 5654
rect 4538 5620 4562 5654
rect 4600 5620 4606 5654
rect 4606 5620 4634 5654
rect 4672 5620 4674 5654
rect 4674 5620 4706 5654
rect 4744 5620 4776 5654
rect 4776 5620 4778 5654
rect 4816 5620 4844 5654
rect 4844 5620 4850 5654
rect 4888 5620 4912 5654
rect 4912 5620 4922 5654
rect 4960 5620 4980 5654
rect 4980 5620 4994 5654
rect 5032 5620 5048 5654
rect 5048 5620 5066 5654
rect 5104 5620 5116 5654
rect 5116 5620 5138 5654
rect 5176 5620 5184 5654
rect 5184 5620 5210 5654
rect 5248 5620 5252 5654
rect 5252 5620 5282 5654
rect 5320 5620 5354 5654
rect 5392 5620 5422 5654
rect 5422 5620 5426 5654
rect 5464 5620 5490 5654
rect 5490 5620 5498 5654
rect 5536 5620 5558 5654
rect 5558 5620 5570 5654
rect 5608 5620 5626 5654
rect 5626 5620 5642 5654
rect 5680 5620 5694 5654
rect 5694 5620 5714 5654
rect 5752 5620 5762 5654
rect 5762 5620 5786 5654
rect 5824 5620 5830 5654
rect 5830 5620 5858 5654
rect 5896 5620 5898 5654
rect 5898 5620 5930 5654
rect 5968 5620 6000 5654
rect 6000 5620 6002 5654
rect 6040 5620 6068 5654
rect 6068 5620 6074 5654
rect 6112 5620 6136 5654
rect 6136 5620 6146 5654
rect 6184 5620 6218 5654
rect 5336 5547 5348 5581
rect 5348 5547 5370 5581
rect 5408 5547 5416 5581
rect 5416 5547 5442 5581
rect 5480 5547 5484 5581
rect 5484 5547 5514 5581
rect 5552 5547 5586 5581
rect 5624 5547 5654 5581
rect 5654 5547 5658 5581
rect 5696 5547 5722 5581
rect 5722 5547 5730 5581
rect 5768 5547 5790 5581
rect 5790 5547 5802 5581
rect 5840 5547 5858 5581
rect 5858 5547 5874 5581
rect 5912 5547 5926 5581
rect 5926 5547 5946 5581
rect 5984 5547 5994 5581
rect 5994 5547 6018 5581
rect 6056 5547 6062 5581
rect 6062 5547 6090 5581
rect 6128 5547 6130 5581
rect 6130 5547 6162 5581
rect 6200 5547 6234 5581
rect 4150 5443 4184 5469
rect 4150 5435 4184 5443
rect 4150 5375 4184 5397
rect 4150 5363 4184 5375
rect 4199 5283 4233 5317
rect 4271 5283 4305 5317
rect 3974 5138 4008 5172
rect 4046 5138 4080 5172
rect 4150 4705 4184 4737
rect 4150 4703 4184 4705
rect 4150 4637 4184 4665
rect 4150 4631 4184 4637
rect 4362 5215 4396 5249
rect 4434 5247 4468 5249
rect 4434 5215 4447 5247
rect 4447 5215 4468 5247
rect 4429 4802 4463 4836
rect 4501 4807 4535 4836
rect 4501 4802 4502 4807
rect 4502 4802 4535 4807
rect 4570 5138 4604 5172
rect 4642 5138 4676 5172
rect 4854 5443 4888 5469
rect 4854 5435 4888 5443
rect 4854 5375 4888 5397
rect 4854 5363 4888 5375
rect 5336 5473 5348 5507
rect 5348 5473 5370 5507
rect 5408 5473 5416 5507
rect 5416 5473 5442 5507
rect 5480 5473 5484 5507
rect 5484 5473 5514 5507
rect 5552 5473 5586 5507
rect 5624 5473 5654 5507
rect 5654 5473 5658 5507
rect 5696 5473 5722 5507
rect 5722 5473 5730 5507
rect 5768 5473 5790 5507
rect 5790 5473 5802 5507
rect 5840 5473 5858 5507
rect 5858 5473 5874 5507
rect 5912 5473 5926 5507
rect 5926 5473 5946 5507
rect 5984 5473 5994 5507
rect 5994 5473 6018 5507
rect 6056 5473 6062 5507
rect 6062 5473 6090 5507
rect 6128 5473 6130 5507
rect 6130 5473 6162 5507
rect 6200 5473 6234 5507
rect 4958 5215 4992 5249
rect 5030 5215 5064 5249
rect 5348 5371 5382 5405
rect 5348 5322 5382 5333
rect 5348 5299 5382 5322
rect 4766 4943 4800 4977
rect 4766 4871 4800 4905
rect 4854 4705 4888 4737
rect 4854 4703 4888 4705
rect 4854 4637 4888 4665
rect 4854 4631 4888 4637
rect 5435 5011 5469 5045
rect 5435 4939 5469 4973
rect 5648 5371 5682 5405
rect 5648 5322 5682 5333
rect 5648 5299 5682 5322
rect 5524 5122 5558 5156
rect 5524 5050 5558 5084
rect 5348 4628 5382 4654
rect 5348 4620 5382 4628
rect 5348 4548 5382 4582
rect 5725 5007 5759 5041
rect 5725 4935 5759 4969
rect 6000 5371 6034 5405
rect 6000 5322 6034 5333
rect 6000 5299 6034 5322
rect 6088 5194 6122 5204
rect 6088 5170 6089 5194
rect 6089 5170 6122 5194
rect 6088 5126 6122 5132
rect 6088 5098 6089 5126
rect 6089 5098 6122 5126
rect 5919 5007 5953 5041
rect 5919 4935 5953 4969
rect 5823 4800 5857 4834
rect 5823 4730 5824 4762
rect 5824 4730 5857 4762
rect 5823 4728 5857 4730
rect 5648 4628 5682 4654
rect 5648 4620 5682 4628
rect 5648 4548 5682 4582
rect 6000 4628 6034 4654
rect 6000 4620 6034 4628
rect 6000 4548 6034 4582
rect 6177 5026 6211 5041
rect 6177 5007 6210 5026
rect 6210 5007 6211 5026
rect 6177 4958 6211 4969
rect 6177 4935 6210 4958
rect 6210 4935 6211 4958
rect 4055 4436 4069 4470
rect 4069 4436 4089 4470
rect 4127 4436 4137 4470
rect 4137 4436 4161 4470
rect 4199 4436 4205 4470
rect 4205 4436 4233 4470
rect 4271 4436 4273 4470
rect 4273 4436 4305 4470
rect 4343 4436 4375 4470
rect 4375 4436 4377 4470
rect 4415 4436 4443 4470
rect 4443 4436 4449 4470
rect 4487 4436 4511 4470
rect 4511 4436 4521 4470
rect 4559 4436 4579 4470
rect 4579 4436 4593 4470
rect 4631 4436 4647 4470
rect 4647 4436 4665 4470
rect 4703 4436 4715 4470
rect 4715 4436 4737 4470
rect 4775 4436 4783 4470
rect 4783 4436 4809 4470
rect 4847 4436 4851 4470
rect 4851 4436 4881 4470
rect 4919 4436 4953 4470
rect 4991 4436 5021 4470
rect 5021 4436 5025 4470
rect 5063 4436 5089 4470
rect 5089 4436 5097 4470
rect 5135 4436 5157 4470
rect 5157 4436 5169 4470
rect 5230 4467 5264 4501
rect 5302 4467 5332 4501
rect 5332 4467 5336 4501
rect 5374 4467 5400 4501
rect 5400 4467 5408 4501
rect 5446 4467 5468 4501
rect 5468 4467 5480 4501
rect 5518 4467 5536 4501
rect 5536 4467 5552 4501
rect 5590 4467 5604 4501
rect 5604 4467 5624 4501
rect 5662 4467 5672 4501
rect 5672 4467 5696 4501
rect 5734 4467 5740 4501
rect 5740 4467 5768 4501
rect 5806 4467 5808 4501
rect 5808 4467 5840 4501
rect 5878 4467 5910 4501
rect 5910 4467 5912 4501
rect 5950 4467 5978 4501
rect 5978 4467 5984 4501
rect 6022 4467 6046 4501
rect 6046 4467 6056 4501
rect 6094 4467 6114 4501
rect 6114 4467 6128 4501
rect 4117 4266 4151 4272
rect 4117 4238 4151 4266
rect 4117 4198 4151 4200
rect 4117 4166 4151 4198
rect 4199 3922 4233 3956
rect 4199 3850 4233 3884
rect 3941 3731 3975 3765
rect 4013 3731 4047 3765
rect 4117 3528 4151 3540
rect 4117 3506 4151 3528
rect 4117 3460 4151 3468
rect 4117 3434 4151 3460
rect 4395 3935 4429 3969
rect 4467 3964 4469 3969
rect 4469 3964 4501 3969
rect 4467 3935 4501 3964
rect 4329 3654 4363 3688
rect 4401 3656 4414 3688
rect 4414 3656 4435 3688
rect 4401 3654 4435 3656
rect 4736 3835 4770 3869
rect 4821 4266 4855 4272
rect 4821 4238 4855 4266
rect 4821 4198 4855 4200
rect 4821 4166 4855 4198
rect 5323 4238 5357 4246
rect 5323 4212 5357 4238
rect 5323 4140 5357 4174
rect 5675 4386 5709 4420
rect 5675 4340 5709 4348
rect 5675 4314 5709 4340
rect 5752 3999 5786 4033
rect 5752 3927 5786 3961
rect 5409 3876 5443 3877
rect 4537 3731 4571 3765
rect 4609 3731 4643 3765
rect 4736 3763 4770 3797
rect 5409 3843 5443 3876
rect 5409 3774 5443 3805
rect 5409 3771 5443 3774
rect 4925 3654 4959 3688
rect 4997 3654 5031 3688
rect 4821 3528 4855 3540
rect 4821 3506 4855 3528
rect 4821 3460 4855 3468
rect 4821 3434 4855 3460
rect 5323 3646 5357 3669
rect 5323 3635 5357 3646
rect 5323 3563 5357 3597
rect 6027 4386 6061 4420
rect 6027 4340 6061 4348
rect 6027 4314 6061 4340
rect 5588 3842 5621 3876
rect 5621 3842 5622 3876
rect 5588 3774 5621 3804
rect 5621 3774 5622 3804
rect 5850 3851 5884 3885
rect 5850 3779 5884 3813
rect 5588 3770 5622 3774
rect 5675 3646 5709 3669
rect 5675 3635 5709 3646
rect 5675 3563 5709 3597
rect 5946 3997 5980 4031
rect 5946 3925 5980 3959
rect 6116 4212 6150 4246
rect 6116 4140 6150 4174
rect 6204 4010 6237 4031
rect 6237 4010 6238 4031
rect 6204 3997 6238 4010
rect 6204 3942 6237 3959
rect 6237 3942 6238 3959
rect 6204 3925 6238 3942
rect 6027 3646 6061 3669
rect 6027 3635 6061 3646
rect 6027 3563 6061 3597
rect 5126 3478 5138 3512
rect 5138 3478 5160 3512
rect 5198 3478 5206 3512
rect 5206 3478 5232 3512
rect 5270 3478 5274 3512
rect 5274 3478 5304 3512
rect 5342 3478 5376 3512
rect 5414 3478 5444 3512
rect 5444 3478 5448 3512
rect 5486 3478 5512 3512
rect 5512 3478 5520 3512
rect 5558 3478 5580 3512
rect 5580 3478 5592 3512
rect 5630 3478 5648 3512
rect 5648 3478 5664 3512
rect 5702 3478 5716 3512
rect 5716 3478 5736 3512
rect 5774 3478 5784 3512
rect 5784 3478 5808 3512
rect 5846 3478 5852 3512
rect 5852 3478 5880 3512
rect 5918 3478 5920 3512
rect 5920 3478 5952 3512
rect 5990 3478 6022 3512
rect 6022 3478 6024 3512
rect 6062 3478 6090 3512
rect 6090 3478 6096 3512
rect 6134 3478 6158 3512
rect 6158 3478 6168 3512
rect 6206 3478 6240 3512
rect -8920 2846 -8886 2880
rect -8920 2800 -8886 2808
rect -8920 2774 -8886 2800
rect -9006 2453 -8972 2487
rect -9180 2336 -9146 2343
rect -9180 2309 -9152 2336
rect -9152 2309 -9146 2336
rect -9180 2268 -9146 2271
rect -9180 2237 -9152 2268
rect -9152 2237 -9146 2268
rect -9096 2302 -9062 2336
rect -9096 2230 -9062 2264
rect -9006 2381 -8972 2415
rect -8744 2504 -8710 2533
rect -8744 2499 -8710 2504
rect -8827 2453 -8793 2487
rect -8827 2381 -8793 2415
rect -8744 2436 -8710 2461
rect -8744 2427 -8710 2436
rect -9272 2106 -9238 2129
rect -9272 2095 -9238 2106
rect -9272 2023 -9238 2057
rect -8568 2846 -8534 2880
rect -8568 2800 -8534 2808
rect -8568 2774 -8534 2800
rect -8649 2302 -8624 2336
rect -8624 2302 -8615 2336
rect -8649 2234 -8624 2264
rect -8624 2234 -8615 2264
rect -8649 2230 -8615 2234
rect -8920 2106 -8886 2129
rect -8920 2095 -8886 2106
rect -8920 2023 -8886 2057
<< metal1 >>
rect 3836 7623 6233 7628
rect 3836 7616 5099 7623
rect 3836 7582 3883 7616
rect 3917 7582 3955 7616
rect 3989 7582 4027 7616
rect 4061 7582 4099 7616
rect 4133 7582 4171 7616
rect 4205 7582 4243 7616
rect 4277 7582 4315 7616
rect 4349 7582 4387 7616
rect 4421 7582 4459 7616
rect 4493 7582 4531 7616
rect 4565 7582 4603 7616
rect 4637 7582 4675 7616
rect 4709 7582 4747 7616
rect 4781 7582 4819 7616
rect 4853 7582 4891 7616
rect 4925 7582 4963 7616
rect 4997 7582 5035 7616
rect 5069 7582 5099 7616
rect 3836 7571 5099 7582
rect 5151 7571 5178 7623
rect 5230 7616 5256 7623
rect 5308 7616 6233 7623
rect 5230 7582 5251 7616
rect 5308 7582 5323 7616
rect 5357 7582 5395 7616
rect 5429 7582 5467 7616
rect 5501 7582 5539 7616
rect 5573 7582 5611 7616
rect 5645 7582 5683 7616
rect 5717 7582 5755 7616
rect 5789 7582 5827 7616
rect 5861 7582 5899 7616
rect 5933 7582 5971 7616
rect 6005 7582 6043 7616
rect 6077 7582 6115 7616
rect 6149 7582 6187 7616
rect 6221 7582 6233 7616
rect 5230 7571 5256 7582
rect 5308 7571 6233 7582
rect 3836 7544 6233 7571
rect 3836 7531 5099 7544
rect 3836 7497 4231 7531
rect 4265 7497 4707 7531
rect 4741 7497 5099 7531
rect 3836 7492 5099 7497
rect 5151 7492 5178 7544
rect 5230 7492 5256 7544
rect 5308 7531 6233 7544
rect 5308 7497 5535 7531
rect 5569 7497 5835 7531
rect 5869 7497 6187 7531
rect 6221 7497 6233 7531
rect 5308 7492 6233 7497
rect 3836 7465 6233 7492
rect 3836 7459 5099 7465
rect 3836 7425 4231 7459
rect 4265 7425 4707 7459
rect 4741 7425 5099 7459
rect 3836 7413 5099 7425
rect 5151 7413 5178 7465
rect 5230 7413 5256 7465
rect 5308 7459 6233 7465
rect 5308 7425 5535 7459
rect 5569 7425 5835 7459
rect 5869 7425 6187 7459
rect 6221 7425 6233 7459
rect 5308 7413 6233 7425
rect 3836 7412 6233 7413
rect 3965 7302 4011 7314
rect 3965 7268 3971 7302
rect 4005 7268 4011 7302
rect 3965 7230 4011 7268
rect 3965 7196 3971 7230
rect 4005 7196 4011 7230
rect 3965 7184 4011 7196
rect 4434 7312 4486 7318
rect 4434 7245 4486 7260
rect 4434 7187 4486 7193
rect 4603 7312 4655 7318
rect 4603 7245 4655 7260
rect 4603 7187 4655 7193
rect 4786 7316 4838 7322
rect 4786 7249 4838 7264
rect 4786 7191 4838 7197
rect 4959 7316 5011 7322
rect 4959 7249 5011 7264
rect 4959 7191 5011 7197
rect 5436 7316 5488 7322
rect 5436 7249 5488 7264
rect 5436 7191 5488 7197
rect 5579 7246 5659 7298
rect 5711 7246 5723 7298
rect 5775 7246 5781 7298
tri 5575 7187 5579 7191 se
rect 5579 7187 5613 7246
tri 5613 7212 5647 7246 nw
tri 5572 7184 5575 7187 se
rect 5575 7184 5613 7187
tri 5567 7179 5572 7184 se
rect 5572 7179 5613 7184
tri 5557 7169 5567 7179 se
rect 5567 7169 5613 7179
rect 4524 7167 4570 7169
tri 4570 7167 4572 7169 sw
tri 5555 7167 5557 7169 se
rect 5557 7167 5613 7169
rect 4524 7157 4572 7167
tri 4572 7157 4582 7167 sw
tri 5545 7157 5555 7167 se
rect 5555 7157 5613 7167
rect 4524 7123 4530 7157
rect 4564 7123 5613 7157
rect 5653 7167 5699 7179
tri 5699 7167 5706 7174 sw
tri 5904 7167 5911 7174 se
rect 5911 7167 5957 7179
tri 5957 7167 5964 7174 sw
tri 6098 7167 6105 7174 se
rect 6105 7167 6151 7179
rect 5653 7133 5659 7167
rect 5693 7140 5706 7167
tri 5706 7140 5733 7167 sw
tri 5877 7140 5904 7167 se
rect 5904 7140 5917 7167
rect 5693 7133 5917 7140
rect 5951 7140 5964 7167
tri 5964 7140 5991 7167 sw
tri 6071 7140 6098 7167 se
rect 6098 7140 6111 7167
rect 5951 7133 6111 7140
rect 6145 7133 6151 7167
rect 4524 7095 4576 7123
tri 4576 7095 4604 7123 nw
rect 5653 7095 6151 7133
rect 4524 7085 4570 7095
tri 4570 7089 4576 7095 nw
rect 4049 7054 4095 7066
rect 4049 7020 4055 7054
rect 4089 7039 4095 7054
rect 4524 7051 4530 7085
rect 4564 7051 4570 7085
tri 4095 7039 4106 7050 sw
rect 4524 7039 4570 7051
rect 4794 7067 5442 7095
rect 4794 7061 4856 7067
tri 4856 7061 4862 7067 nw
tri 5412 7061 5418 7067 ne
rect 5418 7061 5442 7067
rect 4794 7045 4840 7061
tri 4840 7045 4856 7061 nw
tri 5418 7045 5434 7061 ne
rect 5434 7045 5442 7061
tri 4792 7043 4794 7045 se
rect 4794 7043 4838 7045
tri 4838 7043 4840 7045 nw
tri 5434 7043 5436 7045 ne
rect 5436 7043 5442 7045
rect 5494 7043 5506 7095
rect 5558 7043 5564 7095
rect 5653 7061 5659 7095
rect 5693 7076 5917 7095
rect 5693 7061 5711 7076
tri 5711 7061 5726 7076 nw
tri 5884 7061 5899 7076 ne
rect 5899 7061 5917 7076
rect 5951 7076 6111 7095
rect 5951 7061 5969 7076
tri 5969 7061 5984 7076 nw
tri 6078 7061 6093 7076 ne
rect 6093 7061 6111 7076
rect 6145 7061 6151 7095
rect 5653 7049 5699 7061
tri 5699 7049 5711 7061 nw
tri 5899 7049 5911 7061 ne
rect 5911 7049 5957 7061
tri 5957 7049 5969 7061 nw
tri 6093 7049 6105 7061 ne
rect 6105 7049 6151 7061
tri 4788 7039 4792 7043 se
rect 4792 7039 4834 7043
tri 4834 7039 4838 7043 nw
rect 4089 7037 4106 7039
tri 4106 7037 4108 7039 sw
tri 4786 7037 4788 7039 se
rect 4788 7037 4832 7039
tri 4832 7037 4834 7039 nw
rect 4089 7034 4108 7037
tri 4108 7034 4111 7037 sw
tri 4783 7034 4786 7037 se
rect 4786 7034 4829 7037
tri 4829 7034 4832 7037 nw
rect 4089 7027 4111 7034
tri 4111 7027 4118 7034 sw
tri 4776 7027 4783 7034 se
rect 4783 7027 4828 7034
tri 4828 7033 4829 7034 nw
rect 4089 7025 4118 7027
tri 4118 7025 4120 7027 sw
tri 4774 7025 4776 7027 se
rect 4776 7025 4828 7027
rect 4089 7020 4120 7025
rect 4049 7016 4120 7020
tri 4120 7016 4129 7025 sw
tri 4765 7016 4774 7025 se
rect 4774 7016 4828 7025
rect 4049 7011 4414 7016
tri 4414 7011 4419 7016 sw
tri 4760 7011 4765 7016 se
rect 4765 7011 4828 7016
rect 4049 6982 4828 7011
rect 4049 6948 4055 6982
rect 4089 6962 4107 6982
tri 4107 6962 4127 6982 nw
tri 4358 6977 4363 6982 ne
rect 4363 6977 4828 6982
rect 4877 7025 5307 7037
rect 4877 6991 4883 7025
rect 4917 6992 5267 7025
rect 4917 6991 4957 6992
tri 4957 6991 4958 6992 nw
tri 5226 6991 5227 6992 ne
rect 5227 6991 5267 6992
rect 5301 6991 5307 7025
rect 4877 6982 4948 6991
tri 4948 6982 4957 6991 nw
tri 5227 6982 5236 6991 ne
rect 5236 6982 5307 6991
rect 4877 6962 4928 6982
tri 4928 6962 4948 6982 nw
tri 5236 6964 5254 6982 ne
rect 5254 6964 5307 6982
rect 4089 6955 4100 6962
tri 4100 6955 4107 6962 nw
rect 4089 6953 4098 6955
tri 4098 6953 4100 6955 nw
rect 4877 6953 4923 6962
tri 4923 6957 4928 6962 nw
rect 5002 6958 5054 6964
tri 5254 6962 5256 6964 ne
rect 5256 6962 5307 6964
rect 4089 6951 4096 6953
tri 4096 6951 4098 6953 nw
rect 4089 6948 4095 6951
tri 4095 6950 4096 6951 nw
rect 4049 6936 4095 6948
rect 4138 6939 4184 6951
rect 4138 6905 4144 6939
rect 4178 6910 4184 6939
rect 4877 6919 4883 6953
rect 4917 6919 4923 6953
tri 4184 6910 4187 6913 sw
rect 4178 6907 4187 6910
tri 4187 6907 4190 6910 sw
rect 4877 6907 4923 6919
tri 4999 6910 5002 6913 se
tri 4996 6907 4999 6910 se
rect 4999 6907 5002 6910
rect 4178 6905 4190 6907
rect 4138 6879 4190 6905
tri 4190 6879 4218 6907 sw
tri 4968 6879 4996 6907 se
rect 4996 6906 5002 6907
tri 5256 6957 5261 6962 ne
rect 5261 6953 5307 6962
rect 5261 6919 5267 6953
rect 5301 6919 5307 6953
rect 5261 6907 5307 6919
rect 5353 7034 5399 7039
tri 5399 7034 5403 7038 sw
tri 5733 7034 5737 7038 se
rect 5737 7034 5783 7046
rect 5353 7027 5403 7034
rect 5353 6993 5359 7027
rect 5393 7004 5403 7027
tri 5403 7004 5433 7034 sw
tri 5703 7004 5733 7034 se
rect 5733 7004 5743 7034
rect 5393 7000 5743 7004
rect 5777 7000 5783 7034
rect 5393 6993 5783 7000
rect 5353 6962 5783 6993
rect 5353 6958 5743 6962
rect 5353 6955 5403 6958
rect 5353 6921 5359 6955
rect 5393 6928 5403 6955
tri 5403 6928 5433 6958 nw
tri 5695 6928 5725 6958 ne
rect 5725 6928 5743 6958
rect 5777 6928 5783 6962
rect 5393 6921 5399 6928
tri 5399 6924 5403 6928 nw
tri 5725 6924 5729 6928 ne
rect 5729 6924 5783 6928
rect 5353 6909 5399 6921
tri 5729 6916 5737 6924 ne
rect 5737 6916 5783 6924
rect 6005 6982 6051 6994
rect 6005 6948 6011 6982
rect 6045 6948 6051 6982
rect 6005 6910 6051 6948
rect 4996 6894 5054 6906
rect 4996 6879 5002 6894
rect 4138 6867 5002 6879
rect 4138 6833 4144 6867
rect 4178 6842 5002 6867
rect 6005 6876 6011 6910
rect 6045 6876 6051 6910
rect 6005 6864 6051 6876
rect 4178 6836 5054 6842
rect 4178 6833 4184 6836
rect 4138 6821 4184 6833
tri 4184 6821 4199 6836 nw
rect 3836 6780 6233 6793
rect 3836 6746 3879 6780
rect 3913 6746 4231 6780
rect 4265 6746 4355 6780
rect 4389 6746 4707 6780
rect 4741 6746 5059 6780
rect 5093 6746 5183 6780
rect 5217 6746 5535 6780
rect 5569 6746 5835 6780
rect 5869 6746 6187 6780
rect 6221 6746 6233 6780
rect 3836 6708 6233 6746
rect 3836 6674 3879 6708
rect 3913 6674 4231 6708
rect 4265 6674 4355 6708
rect 4389 6674 4707 6708
rect 4741 6674 5059 6708
rect 5093 6674 5183 6708
rect 5217 6674 5535 6708
rect 5569 6674 5835 6708
rect 5869 6674 6187 6708
rect 6221 6674 6233 6708
rect 3836 6635 6233 6674
rect 3836 6601 3883 6635
rect 3917 6601 3955 6635
rect 3989 6601 4027 6635
rect 4061 6601 4099 6635
rect 4133 6601 4171 6635
rect 4205 6601 4243 6635
rect 4277 6601 4315 6635
rect 4349 6601 4387 6635
rect 4421 6601 4459 6635
rect 4493 6601 4531 6635
rect 4565 6601 4603 6635
rect 4637 6601 4675 6635
rect 4709 6601 4747 6635
rect 4781 6601 4819 6635
rect 4853 6601 4891 6635
rect 4925 6601 4963 6635
rect 4997 6601 5035 6635
rect 5069 6601 5107 6635
rect 5141 6601 5179 6635
rect 5213 6601 5251 6635
rect 5285 6601 5323 6635
rect 5357 6601 5395 6635
rect 5429 6601 5467 6635
rect 5501 6601 5539 6635
rect 5573 6601 5611 6635
rect 5645 6601 5683 6635
rect 5717 6601 5755 6635
rect 5789 6601 5827 6635
rect 5861 6601 5899 6635
rect 5933 6601 5971 6635
rect 6005 6601 6043 6635
rect 6077 6601 6115 6635
rect 6149 6601 6233 6635
rect 3836 6590 6233 6601
tri 3836 6562 3864 6590 ne
rect 3864 6562 6233 6590
tri 3864 6559 3867 6562 ne
rect 3867 6528 4231 6562
rect 4265 6528 4355 6562
rect 4389 6528 4707 6562
rect 4741 6528 4831 6562
rect 4865 6528 5183 6562
rect 5217 6528 5535 6562
rect 5569 6528 5835 6562
rect 5869 6528 6187 6562
rect 6221 6528 6233 6562
rect 3867 6490 6233 6528
rect 3867 6456 4231 6490
rect 4265 6456 4355 6490
rect 4389 6456 4707 6490
rect 4741 6456 4831 6490
rect 4865 6456 5183 6490
rect 5217 6456 5535 6490
rect 5569 6456 5835 6490
rect 5869 6456 6187 6490
rect 6221 6456 6233 6490
rect 3867 6443 6233 6456
rect 6005 6380 6051 6392
rect 4134 6346 4180 6349
tri 4180 6346 4183 6349 sw
rect 6005 6346 6011 6380
rect 6045 6346 6051 6380
rect 4134 6340 4183 6346
tri 4183 6340 4189 6346 sw
tri 5266 6340 5268 6342 se
rect 5268 6340 5314 6342
rect 4134 6337 4564 6340
rect 4134 6303 4140 6337
rect 4174 6303 4564 6337
tri 5262 6336 5266 6340 se
rect 5266 6336 5314 6340
rect 4134 6294 4564 6303
rect 4134 6274 4194 6294
tri 4194 6274 4214 6294 nw
tri 4484 6274 4504 6294 ne
rect 4504 6274 4564 6294
rect 4134 6265 4182 6274
rect 4134 6231 4140 6265
rect 4174 6262 4182 6265
tri 4182 6262 4194 6274 nw
tri 4504 6262 4516 6274 ne
rect 4516 6262 4564 6274
rect 4174 6231 4180 6262
tri 4180 6260 4182 6262 nw
tri 4516 6260 4518 6262 ne
rect 4134 6219 4180 6231
rect 4433 6246 4479 6258
rect 4433 6212 4439 6246
rect 4473 6212 4479 6246
tri 4412 6187 4433 6208 se
rect 4433 6187 4479 6212
tri 4400 6175 4412 6187 se
rect 4412 6175 4479 6187
tri 4399 6174 4400 6175 se
rect 4400 6174 4479 6175
rect 4049 6140 4439 6174
rect 4473 6140 4479 6174
rect 4049 6128 4479 6140
rect 4518 6208 4564 6262
rect 4695 6330 5314 6336
rect 4747 6296 5274 6330
rect 5308 6296 5314 6330
rect 4747 6284 5314 6296
rect 4747 6278 4771 6284
rect 4695 6274 4771 6278
tri 4771 6274 4781 6284 nw
tri 5234 6274 5244 6284 ne
rect 5244 6274 5314 6284
rect 4695 6266 4759 6274
rect 4747 6262 4759 6266
tri 4759 6262 4771 6274 nw
tri 5244 6262 5256 6274 ne
rect 5256 6262 5314 6274
rect 6005 6308 6051 6346
rect 6005 6274 6011 6308
rect 6045 6274 6051 6308
rect 6005 6262 6051 6274
rect 4747 6258 4755 6262
tri 4755 6258 4759 6262 nw
tri 5256 6258 5260 6262 ne
rect 5260 6258 5314 6262
tri 4747 6250 4755 6258 nw
tri 5260 6250 5268 6258 ne
tri 4564 6208 4570 6214 sw
rect 4695 6208 4747 6214
rect 4786 6240 4838 6246
rect 4518 6206 4570 6208
tri 4570 6206 4572 6208 sw
rect 4518 6187 4572 6206
tri 4572 6187 4591 6206 sw
tri 4767 6187 4786 6206 se
rect 4786 6187 4838 6188
rect 4518 6180 4591 6187
tri 4591 6180 4598 6187 sw
tri 4760 6180 4767 6187 se
rect 4767 6180 4838 6187
rect 4518 6176 4838 6180
rect 4518 6134 4786 6176
tri 4770 6128 4776 6134 ne
rect 4776 6128 4786 6134
rect 4049 6115 4116 6128
tri 4116 6115 4129 6128 nw
tri 4776 6118 4786 6128 ne
rect 4786 6118 4838 6124
rect 5001 6227 5054 6233
rect 5001 6175 5002 6227
rect 5268 6224 5274 6258
rect 5308 6224 5314 6258
rect 5268 6212 5314 6224
rect 5001 6161 5054 6175
rect 4049 6109 4110 6115
tri 4110 6109 4116 6115 nw
rect 5001 6109 5002 6161
rect 5653 6175 5699 6187
tri 5699 6175 5711 6187 sw
tri 5899 6175 5911 6187 se
rect 5911 6175 5957 6187
tri 5957 6175 5969 6187 sw
tri 6093 6175 6105 6187 se
rect 6105 6175 6151 6187
rect 4049 6103 4104 6109
tri 4104 6103 4110 6109 nw
rect 5001 6103 5054 6109
rect 5087 6143 5133 6155
tri 5133 6143 5137 6147 sw
tri 5349 6143 5353 6147 se
rect 5353 6143 5399 6155
rect 5087 6109 5093 6143
rect 5127 6113 5137 6143
tri 5137 6113 5167 6143 sw
tri 5319 6113 5349 6143 se
rect 5349 6113 5359 6143
rect 5127 6109 5359 6113
rect 5393 6109 5399 6143
rect 4049 6102 4095 6103
rect 4049 6068 4055 6102
rect 4089 6068 4095 6102
tri 4095 6094 4104 6103 nw
rect 4049 6030 4095 6068
rect 3956 6017 4002 6029
rect 3956 5983 3962 6017
rect 3996 5983 4002 6017
rect 4049 5996 4055 6030
rect 4089 5996 4095 6030
rect 4049 5984 4095 5996
rect 4176 6030 4821 6076
rect 4176 6022 4261 6030
tri 4261 6022 4269 6030 nw
tri 4791 6024 4797 6030 ne
rect 4797 6024 4821 6030
rect 4873 6024 4885 6076
rect 4937 6024 4943 6076
rect 5087 6071 5399 6109
rect 5087 6037 5093 6071
rect 5127 6067 5359 6071
rect 5127 6037 5137 6067
tri 5137 6037 5167 6067 nw
tri 5319 6037 5349 6067 ne
rect 5349 6037 5359 6067
rect 5393 6037 5399 6071
rect 5653 6141 5659 6175
rect 5693 6160 5711 6175
tri 5711 6160 5726 6175 sw
tri 5884 6160 5899 6175 se
rect 5899 6160 5917 6175
rect 5693 6141 5917 6160
rect 5951 6160 5969 6175
tri 5969 6160 5984 6175 sw
tri 6078 6160 6093 6175 se
rect 6093 6160 6111 6175
rect 5951 6141 6111 6160
rect 6145 6141 6151 6175
rect 5653 6103 6151 6141
rect 5653 6069 5659 6103
rect 5693 6096 5917 6103
rect 5693 6069 5706 6096
tri 5706 6069 5733 6096 nw
tri 5877 6069 5904 6096 ne
rect 5904 6069 5917 6096
rect 5951 6096 6111 6103
rect 5951 6069 5964 6096
tri 5964 6069 5991 6096 nw
tri 6071 6069 6098 6096 ne
rect 6098 6069 6111 6096
rect 6145 6069 6151 6103
rect 5653 6057 5699 6069
tri 5699 6062 5706 6069 nw
tri 5904 6062 5911 6069 ne
rect 5911 6057 5957 6069
tri 5957 6062 5964 6069 nw
tri 6098 6062 6105 6069 ne
rect 6105 6057 6151 6069
rect 5087 6025 5133 6037
tri 5133 6033 5137 6037 nw
tri 5349 6033 5353 6037 ne
rect 5353 6025 5399 6037
rect 5729 6033 5781 6039
rect 4176 5997 4236 6022
tri 4236 5997 4261 6022 nw
rect 3956 5951 4002 5983
tri 4002 5951 4030 5979 sw
tri 4148 5951 4176 5979 se
rect 4176 5951 4235 5997
tri 4235 5996 4236 5997 nw
rect 3956 5950 4030 5951
tri 4030 5950 4031 5951 sw
tri 4147 5950 4148 5951 se
rect 4148 5950 4235 5951
rect 3956 5945 4031 5950
tri 4031 5945 4036 5950 sw
tri 4142 5945 4147 5950 se
rect 4147 5945 4235 5950
rect 3956 5911 3962 5945
rect 3996 5911 4235 5945
rect 3956 5899 4235 5911
rect 4519 5991 4655 5997
rect 4571 5985 4655 5991
rect 4571 5951 4615 5985
rect 4649 5951 4655 5985
rect 4571 5939 4655 5951
rect 4695 5990 4983 5996
rect 4695 5956 4707 5990
rect 4741 5956 4779 5990
rect 4813 5956 4865 5990
rect 4899 5956 4937 5990
rect 4971 5956 4983 5990
rect 5440 5993 5572 5999
rect 5440 5987 5520 5993
rect 5356 5976 5408 5982
rect 4695 5950 4983 5956
tri 5347 5953 5356 5962 se
tri 5344 5950 5347 5953 se
rect 5347 5950 5356 5953
rect 4519 5925 4655 5939
rect 4571 5922 4655 5925
tri 4655 5922 4683 5950 sw
tri 5316 5922 5344 5950 se
rect 5344 5924 5356 5950
rect 5344 5922 5408 5924
rect 4571 5913 5408 5922
rect 4571 5879 4615 5913
rect 4649 5912 5408 5913
rect 4649 5879 5356 5912
rect 4571 5876 5356 5879
rect 4571 5873 4659 5876
rect 4519 5871 4659 5873
tri 4659 5871 4664 5876 nw
tri 5334 5871 5339 5876 ne
rect 5339 5871 5356 5876
rect 4519 5867 4655 5871
tri 4655 5867 4659 5871 nw
tri 5339 5867 5343 5871 ne
rect 5343 5867 5356 5871
tri 5343 5854 5356 5867 ne
rect 5440 5953 5446 5987
rect 5480 5953 5520 5987
rect 5440 5941 5520 5953
rect 5440 5929 5572 5941
rect 5440 5915 5520 5929
rect 5440 5881 5446 5915
rect 5480 5881 5520 5915
rect 5440 5877 5520 5881
rect 5729 5962 5781 5981
rect 5729 5904 5781 5910
rect 5440 5865 5572 5877
rect 5356 5854 5408 5860
rect 3867 5819 6265 5825
rect 3867 5811 5095 5819
rect 3867 5777 3879 5811
rect 3913 5777 4231 5811
rect 4265 5777 4355 5811
rect 4389 5777 5095 5811
rect 3867 5767 5095 5777
rect 5147 5767 5178 5819
rect 5230 5767 5261 5819
rect 5313 5811 6265 5819
rect 5313 5777 5835 5811
rect 5869 5777 6187 5811
rect 6221 5777 6265 5811
rect 5313 5767 6265 5777
rect 3867 5753 6265 5767
rect 3867 5739 5095 5753
rect 3867 5705 3879 5739
rect 3913 5705 4231 5739
rect 4265 5705 4355 5739
rect 4389 5705 5095 5739
rect 3867 5701 5095 5705
rect 5147 5701 5178 5753
rect 5230 5701 5261 5753
rect 5313 5739 6265 5753
rect 5313 5705 5835 5739
rect 5869 5705 6187 5739
rect 6221 5705 6265 5739
rect 5313 5701 6265 5705
rect 3867 5687 6265 5701
rect 3867 5654 5095 5687
rect 5147 5654 5178 5687
rect 5230 5654 5261 5687
rect 5313 5654 6265 5687
rect 3867 5620 3880 5654
rect 3914 5620 3952 5654
rect 3986 5620 4024 5654
rect 4058 5620 4096 5654
rect 4130 5620 4168 5654
rect 4202 5620 4240 5654
rect 4274 5620 4312 5654
rect 4346 5620 4384 5654
rect 4418 5620 4456 5654
rect 4490 5620 4528 5654
rect 4562 5620 4600 5654
rect 4634 5620 4672 5654
rect 4706 5620 4744 5654
rect 4778 5620 4816 5654
rect 4850 5620 4888 5654
rect 4922 5620 4960 5654
rect 4994 5620 5032 5654
rect 5066 5635 5095 5654
rect 5147 5635 5176 5654
rect 5230 5635 5248 5654
rect 5313 5635 5320 5654
rect 5066 5621 5104 5635
rect 5138 5621 5176 5635
rect 5210 5621 5248 5635
rect 5282 5621 5320 5635
rect 5066 5620 5095 5621
rect 5147 5620 5176 5621
rect 5230 5620 5248 5621
rect 5313 5620 5320 5621
rect 5354 5620 5392 5654
rect 5426 5620 5464 5654
rect 5498 5620 5536 5654
rect 5570 5620 5608 5654
rect 5642 5620 5680 5654
rect 5714 5620 5752 5654
rect 5786 5620 5824 5654
rect 5858 5620 5896 5654
rect 5930 5620 5968 5654
rect 6002 5620 6040 5654
rect 6074 5620 6112 5654
rect 6146 5620 6184 5654
rect 6218 5620 6265 5654
rect 3867 5569 5095 5620
rect 5147 5569 5178 5620
rect 5230 5569 5261 5620
rect 5313 5581 6265 5620
rect 5313 5569 5336 5581
rect 3867 5555 5336 5569
rect 3867 5503 5095 5555
rect 5147 5503 5178 5555
rect 5230 5503 5261 5555
rect 5313 5547 5336 5555
rect 5370 5547 5408 5581
rect 5442 5547 5480 5581
rect 5514 5547 5552 5581
rect 5586 5547 5624 5581
rect 5658 5547 5696 5581
rect 5730 5547 5768 5581
rect 5802 5547 5840 5581
rect 5874 5547 5912 5581
rect 5946 5547 5984 5581
rect 6018 5547 6056 5581
rect 6090 5547 6128 5581
rect 6162 5547 6200 5581
rect 6234 5547 6265 5581
rect 5313 5507 6265 5547
rect 5313 5503 5336 5507
rect 3867 5489 5336 5503
rect 3867 5469 5095 5489
rect 3867 5435 4150 5469
rect 4184 5435 4854 5469
rect 4888 5437 5095 5469
rect 5147 5437 5178 5489
rect 5230 5437 5261 5489
rect 5313 5473 5336 5489
rect 5370 5473 5408 5507
rect 5442 5473 5480 5507
rect 5514 5473 5552 5507
rect 5586 5473 5624 5507
rect 5658 5473 5696 5507
rect 5730 5473 5768 5507
rect 5802 5473 5840 5507
rect 5874 5473 5912 5507
rect 5946 5473 5984 5507
rect 6018 5473 6056 5507
rect 6090 5473 6128 5507
rect 6162 5473 6200 5507
rect 6234 5473 6265 5507
rect 5313 5437 6265 5473
rect 4888 5435 6265 5437
rect 3867 5424 6265 5435
rect 3867 5397 5095 5424
rect 3867 5363 4150 5397
rect 4184 5363 4854 5397
rect 4888 5372 5095 5397
rect 5147 5372 5178 5424
rect 5230 5372 5261 5424
rect 5313 5405 6265 5424
rect 5313 5372 5348 5405
rect 4888 5371 5348 5372
rect 5382 5371 5648 5405
rect 5682 5371 6000 5405
rect 6034 5371 6265 5405
rect 4888 5363 6265 5371
rect 3867 5351 6265 5363
tri 5218 5333 5236 5351 ne
rect 5236 5333 6265 5351
tri 5236 5323 5246 5333 ne
rect 5246 5323 5348 5333
rect 3816 5271 3822 5323
rect 3874 5271 3886 5323
rect 3938 5317 4317 5323
rect 3938 5283 4199 5317
rect 4233 5283 4271 5317
rect 4305 5283 4317 5317
tri 5246 5299 5270 5323 ne
rect 5270 5299 5348 5323
rect 5382 5299 5648 5333
rect 5682 5299 6000 5333
rect 6034 5299 6265 5333
tri 5270 5287 5282 5299 ne
rect 5282 5287 6265 5299
rect 3938 5277 4317 5283
rect 3938 5271 3962 5277
tri 3962 5271 3968 5277 nw
rect 4350 5249 5076 5255
rect 4350 5215 4362 5249
rect 4396 5215 4434 5249
rect 4468 5215 4958 5249
rect 4992 5215 5030 5249
rect 5064 5215 5076 5249
rect 4350 5209 5076 5215
rect 6082 5204 6128 5216
tri 6076 5178 6082 5184 se
rect 6082 5178 6088 5204
rect 3962 5172 4688 5178
rect 3962 5138 3974 5172
rect 4008 5138 4046 5172
rect 4080 5138 4570 5172
rect 4604 5138 4642 5172
rect 4676 5138 4688 5172
tri 6068 5170 6076 5178 se
rect 6076 5170 6088 5178
rect 6122 5170 6128 5204
tri 6066 5168 6068 5170 se
rect 6068 5168 6128 5170
rect 3962 5132 4688 5138
rect 5518 5156 5564 5168
rect 5518 5122 5524 5156
rect 5558 5154 5564 5156
tri 5564 5154 5578 5168 sw
tri 6052 5154 6066 5168 se
rect 6066 5154 6128 5168
rect 5558 5132 6128 5154
rect 5558 5122 6088 5132
rect 5518 5120 6088 5122
rect 4434 5098 4486 5104
tri 4486 5098 4492 5104 sw
rect 5518 5098 5576 5120
tri 5576 5098 5598 5120 nw
tri 6048 5098 6070 5120 ne
rect 6070 5098 6088 5120
rect 6122 5098 6128 5132
rect 4486 5084 4492 5098
tri 4492 5084 4506 5098 sw
rect 5518 5084 5564 5098
tri 5564 5086 5576 5098 nw
tri 6070 5086 6082 5098 ne
rect 6082 5086 6128 5098
rect 4486 5069 4506 5084
tri 4506 5069 4521 5084 sw
rect 4486 5046 5225 5069
rect 4434 5034 5225 5046
rect 4486 5017 5225 5034
rect 4486 5011 4510 5017
tri 4510 5011 4516 5017 nw
tri 5097 5011 5103 5017 ne
rect 5103 5011 5225 5017
rect 4486 5007 4506 5011
tri 4506 5007 4510 5011 nw
tri 5103 5007 5107 5011 ne
rect 5107 5007 5225 5011
rect 4486 4989 4488 5007
tri 4488 4989 4506 5007 nw
tri 5107 4989 5125 5007 ne
rect 5125 4989 5225 5007
tri 4486 4987 4488 4989 nw
rect 4434 4976 4486 4982
rect 4528 4937 4534 4989
rect 4586 4937 4598 4989
rect 4650 4977 4806 4989
rect 4650 4943 4766 4977
rect 4800 4943 4806 4977
tri 5125 4973 5141 4989 ne
rect 5141 4973 5225 4989
rect 4650 4937 4806 4943
tri 5141 4941 5173 4973 ne
tri 4726 4935 4728 4937 ne
rect 4728 4935 4806 4937
tri 4728 4923 4740 4935 ne
rect 4740 4923 4806 4935
tri 4740 4905 4758 4923 ne
rect 4758 4905 4806 4923
tri 4758 4903 4760 4905 ne
rect 4760 4871 4766 4905
rect 4800 4871 4806 4905
rect 4760 4859 4806 4871
rect 5173 4903 5225 4973
rect 5429 5051 5488 5057
rect 5429 5045 5436 5051
rect 5429 5011 5435 5045
rect 5518 5050 5524 5084
rect 5558 5050 5564 5084
rect 5518 5038 5564 5050
rect 5719 5041 5765 5053
tri 5912 5047 5913 5048 se
rect 5913 5047 5959 5053
tri 5765 5041 5771 5047 sw
tri 5906 5041 5912 5047 se
rect 5912 5041 5959 5047
tri 5959 5041 5966 5048 sw
tri 6164 5041 6171 5048 se
rect 6171 5041 6217 5053
rect 5429 4999 5436 5011
rect 5429 4985 5488 4999
rect 5429 4973 5436 4985
rect 5429 4939 5435 4973
rect 5429 4933 5436 4939
rect 5429 4927 5488 4933
rect 5719 5007 5725 5041
rect 5759 5014 5771 5041
tri 5771 5014 5798 5041 sw
tri 5879 5014 5906 5041 se
rect 5906 5014 5919 5041
rect 5759 5007 5919 5014
rect 5953 5014 5966 5041
tri 5966 5014 5993 5041 sw
tri 6137 5014 6164 5041 se
rect 6164 5014 6177 5041
rect 5953 5007 6177 5014
rect 6211 5007 6217 5041
rect 5719 4969 6217 5007
rect 5719 4935 5725 4969
rect 5759 4950 5919 4969
rect 5759 4935 5777 4950
tri 5777 4935 5792 4950 nw
tri 5886 4935 5901 4950 ne
rect 5901 4935 5919 4950
rect 5953 4950 6177 4969
rect 5953 4935 5971 4950
tri 5971 4935 5986 4950 nw
tri 6144 4935 6159 4950 ne
rect 6159 4935 6177 4950
rect 6211 4935 6217 4969
rect 5719 4923 5765 4935
tri 5765 4923 5777 4935 nw
tri 5901 4923 5913 4935 ne
rect 5913 4923 5959 4935
tri 5959 4923 5971 4935 nw
tri 6159 4923 6171 4935 ne
rect 6171 4923 6217 4935
tri 5225 4903 5239 4917 sw
rect 5520 4912 5572 4918
rect 5173 4869 5239 4903
tri 5239 4869 5273 4903 sw
tri 5486 4869 5520 4903 se
rect 5173 4860 5520 4869
rect 5173 4848 5572 4860
tri 4547 4842 4553 4848 se
rect 4553 4842 4565 4848
rect 4417 4836 4565 4842
rect 4417 4802 4429 4836
rect 4463 4802 4501 4836
rect 4535 4802 4565 4836
rect 4417 4796 4565 4802
rect 4617 4796 4629 4848
rect 4681 4796 4687 4848
rect 5173 4799 5520 4848
tri 5511 4796 5514 4799 ne
rect 5514 4796 5520 4799
tri 5514 4790 5520 4796 ne
rect 5520 4790 5572 4796
rect 5733 4840 5863 4846
rect 5785 4834 5863 4840
rect 5785 4800 5823 4834
rect 5857 4800 5863 4834
rect 5785 4788 5863 4800
rect 5733 4774 5863 4788
tri 4132 4737 4144 4749 se
rect 4144 4737 4894 4749
tri 4098 4703 4132 4737 se
rect 4132 4703 4150 4737
rect 4184 4703 4854 4737
rect 4888 4728 4894 4737
tri 4894 4728 4915 4749 sw
rect 4888 4703 4915 4728
tri 4062 4667 4098 4703 se
rect 4098 4667 4915 4703
tri 4915 4667 4976 4728 sw
rect 5785 4762 5863 4774
rect 5785 4728 5823 4762
rect 5857 4728 5863 4762
rect 5785 4722 5863 4728
rect 5733 4716 5863 4722
tri 4060 4665 4062 4667 se
rect 4062 4665 6292 4667
tri 4044 4649 4060 4665 se
rect 4060 4649 4150 4665
rect 3868 4631 4150 4649
rect 4184 4631 4854 4665
rect 4888 4654 6292 4665
rect 4888 4631 5348 4654
rect 3868 4620 5348 4631
rect 5382 4620 5648 4654
rect 5682 4620 6000 4654
rect 6034 4620 6292 4654
rect 3868 4582 6292 4620
rect 3868 4548 5348 4582
rect 5382 4548 5648 4582
rect 5682 4548 6000 4582
rect 6034 4548 6292 4582
rect 3868 4501 6292 4548
rect 3868 4470 5230 4501
rect 3868 4436 4055 4470
rect 4089 4436 4127 4470
rect 4161 4436 4199 4470
rect 4233 4436 4271 4470
rect 4305 4436 4343 4470
rect 4377 4436 4415 4470
rect 4449 4436 4487 4470
rect 4521 4436 4559 4470
rect 4593 4436 4631 4470
rect 4665 4436 4703 4470
rect 4737 4436 4775 4470
rect 4809 4436 4847 4470
rect 4881 4436 4919 4470
rect 4953 4436 4991 4470
rect 5025 4436 5063 4470
rect 5097 4436 5135 4470
rect 5169 4467 5230 4470
rect 5264 4467 5302 4501
rect 5336 4467 5374 4501
rect 5408 4467 5446 4501
rect 5480 4467 5518 4501
rect 5552 4467 5590 4501
rect 5624 4467 5662 4501
rect 5696 4467 5734 4501
rect 5768 4467 5806 4501
rect 5840 4467 5878 4501
rect 5912 4467 5950 4501
rect 5984 4467 6022 4501
rect 6056 4467 6094 4501
rect 6128 4467 6292 4501
rect 5169 4436 6292 4467
rect 3868 4420 6292 4436
rect 3868 4386 5675 4420
rect 5709 4386 6027 4420
rect 6061 4386 6292 4420
rect 3868 4348 6292 4386
rect 3868 4314 5675 4348
rect 5709 4314 6027 4348
rect 6061 4314 6292 4348
rect 3868 4303 6292 4314
tri 3995 4272 4026 4303 ne
rect 4026 4301 6292 4303
rect 4026 4272 4965 4301
tri 4026 4258 4040 4272 ne
rect 4040 4258 4117 4272
tri 4040 4238 4060 4258 ne
rect 4060 4238 4117 4258
rect 4151 4238 4821 4272
rect 4855 4258 4965 4272
tri 4965 4258 5008 4301 nw
rect 4855 4246 4953 4258
tri 4953 4246 4965 4258 nw
rect 5317 4246 5363 4258
rect 6109 4252 6161 4258
tri 5363 4246 5367 4250 sw
tri 6105 4246 6109 4250 se
rect 4855 4238 4919 4246
tri 4060 4212 4086 4238 ne
rect 4086 4212 4919 4238
tri 4919 4212 4953 4246 nw
rect 5317 4212 5323 4246
rect 5357 4216 5367 4246
tri 5367 4216 5397 4246 sw
tri 6075 4216 6105 4246 se
rect 6105 4216 6109 4246
rect 5357 4212 6109 4216
tri 4086 4200 4098 4212 ne
rect 4098 4200 4881 4212
tri 4098 4187 4111 4200 ne
rect 4111 4166 4117 4200
rect 4151 4166 4821 4200
rect 4855 4174 4881 4200
tri 4881 4174 4919 4212 nw
rect 5317 4200 6109 4212
rect 5317 4183 6161 4200
rect 5317 4174 6109 4183
rect 4855 4166 4861 4174
rect 4111 4154 4861 4166
tri 4861 4154 4881 4174 nw
rect 5317 4140 5323 4174
rect 5357 4170 6109 4174
rect 5357 4140 5367 4170
tri 5367 4140 5397 4170 nw
tri 6075 4140 6105 4170 ne
rect 6105 4140 6109 4170
rect 5317 4128 5363 4140
tri 5363 4136 5367 4140 nw
tri 6105 4136 6109 4140 ne
rect 6109 4125 6161 4131
rect 5746 4033 5792 4045
tri 5939 4042 5940 4043 se
rect 5940 4042 5986 4043
rect 5746 3999 5752 4033
rect 5786 4031 5792 4033
tri 5792 4031 5803 4042 sw
tri 5928 4031 5939 4042 se
rect 5939 4031 5986 4042
tri 5986 4031 5998 4043 sw
tri 6186 4031 6198 4043 se
rect 6198 4031 6244 4043
rect 5786 4016 5803 4031
tri 5803 4016 5818 4031 sw
tri 5913 4016 5928 4031 se
rect 5928 4016 5946 4031
rect 5786 3999 5946 4016
rect 5746 3997 5946 3999
rect 5980 4016 5998 4031
tri 5998 4016 6013 4031 sw
tri 6171 4016 6186 4031 se
rect 6186 4016 6204 4031
rect 5980 3997 6204 4016
rect 6238 3997 6244 4031
rect 4383 3969 5628 3975
rect 3952 3962 4004 3968
tri 4181 3956 4193 3968 se
rect 4193 3956 4239 3968
tri 4172 3947 4181 3956 se
rect 4181 3947 4199 3956
tri 4004 3922 4029 3947 sw
tri 4147 3922 4172 3947 se
rect 4172 3922 4199 3947
rect 4233 3922 4239 3956
rect 4383 3935 4395 3969
rect 4429 3935 4467 3969
rect 4501 3935 5628 3969
rect 4383 3929 5628 3935
tri 5548 3927 5550 3929 ne
rect 5550 3927 5628 3929
tri 5550 3925 5552 3927 ne
rect 5552 3925 5628 3927
rect 4004 3913 4029 3922
tri 4029 3913 4038 3922 sw
tri 4138 3913 4147 3922 se
rect 4147 3913 4239 3922
tri 5552 3915 5562 3925 ne
rect 5562 3915 5628 3925
rect 5746 3961 6244 3997
rect 5746 3927 5752 3961
rect 5786 3959 6244 3961
rect 5786 3952 5946 3959
rect 5786 3927 5799 3952
rect 5746 3925 5799 3927
tri 5799 3925 5826 3952 nw
tri 5901 3925 5928 3952 ne
rect 5928 3925 5946 3952
rect 5980 3952 6204 3959
rect 5980 3925 5998 3952
tri 5998 3925 6025 3952 nw
tri 6165 3925 6192 3952 ne
rect 6192 3925 6204 3952
rect 6238 3925 6244 3959
rect 5746 3915 5792 3925
tri 5792 3918 5799 3925 nw
tri 5928 3918 5935 3925 ne
rect 5935 3918 5986 3925
tri 5935 3915 5938 3918 ne
rect 5938 3915 5986 3918
tri 5562 3913 5564 3915 ne
rect 5564 3913 5628 3915
tri 5938 3913 5940 3915 ne
rect 5940 3913 5986 3915
tri 5986 3913 5998 3925 nw
tri 6192 3919 6198 3925 ne
rect 6198 3913 6244 3925
rect 4004 3910 4239 3913
rect 3952 3898 4239 3910
rect 4004 3884 4239 3898
tri 5564 3897 5580 3913 ne
rect 5580 3897 5628 3913
tri 5580 3895 5582 3897 ne
rect 4004 3861 4199 3884
rect 4004 3850 4014 3861
tri 4014 3850 4025 3861 nw
tri 4170 3850 4181 3861 ne
rect 4181 3850 4199 3861
rect 4233 3850 4239 3884
rect 3952 3840 4004 3846
tri 4004 3840 4014 3850 nw
tri 4181 3840 4191 3850 ne
rect 4191 3840 4239 3850
tri 4191 3838 4193 3840 ne
rect 4193 3838 4239 3840
rect 4358 3829 4364 3881
rect 4416 3829 4428 3881
rect 4480 3869 4776 3881
rect 4480 3835 4736 3869
rect 4770 3835 4776 3869
rect 4480 3829 4776 3835
tri 4696 3813 4712 3829 ne
rect 4712 3813 4776 3829
tri 4712 3805 4720 3813 ne
rect 4720 3805 4776 3813
tri 4720 3797 4728 3805 ne
rect 4728 3797 4776 3805
tri 4728 3795 4730 3797 ne
rect 3929 3765 4655 3771
rect 3929 3731 3941 3765
rect 3975 3731 4013 3765
rect 4047 3731 4537 3765
rect 4571 3731 4609 3765
rect 4643 3731 4655 3765
rect 4730 3763 4736 3797
rect 4770 3763 4776 3797
rect 4730 3751 4776 3763
rect 4891 3877 4943 3882
tri 4943 3877 4947 3881 sw
rect 5403 3877 5449 3889
rect 4891 3876 4947 3877
rect 4943 3871 4947 3876
tri 4947 3871 4953 3877 sw
rect 4943 3843 4953 3871
tri 4953 3843 4981 3871 sw
tri 5375 3843 5403 3871 se
rect 5403 3843 5409 3877
rect 5443 3843 5449 3877
rect 4943 3842 4981 3843
tri 4981 3842 4982 3843 sw
tri 5374 3842 5375 3843 se
rect 5375 3842 5449 3843
rect 4943 3837 4982 3842
tri 4982 3837 4987 3842 sw
tri 5369 3837 5374 3842 se
rect 5374 3837 5449 3842
rect 4943 3824 5449 3837
rect 4891 3812 5449 3824
rect 4943 3805 5449 3812
rect 4943 3799 5409 3805
rect 4943 3795 4964 3799
tri 4964 3795 4968 3799 nw
tri 5369 3795 5373 3799 ne
rect 5373 3795 5409 3799
tri 4943 3774 4964 3795 nw
tri 5373 3774 5394 3795 ne
rect 5394 3774 5409 3795
tri 5394 3771 5397 3774 ne
rect 5397 3771 5409 3774
rect 5443 3771 5449 3805
tri 5397 3770 5398 3771 ne
rect 5398 3770 5449 3771
tri 5398 3765 5403 3770 ne
rect 4891 3754 4943 3760
rect 5403 3759 5449 3770
rect 5582 3876 5628 3897
rect 5582 3842 5588 3876
rect 5622 3842 5628 3876
rect 5582 3804 5628 3842
rect 5582 3770 5588 3804
rect 5622 3770 5628 3804
rect 5582 3758 5628 3770
rect 5814 3891 5890 3897
rect 5866 3885 5890 3891
rect 5884 3851 5890 3885
rect 5866 3839 5890 3851
rect 5814 3825 5890 3839
rect 5866 3813 5890 3825
rect 5884 3779 5890 3813
rect 5866 3773 5890 3779
rect 5814 3767 5890 3773
rect 3929 3725 4655 3731
rect 4317 3688 5043 3694
rect 4317 3654 4329 3688
rect 4363 3654 4401 3688
rect 4435 3654 4925 3688
rect 4959 3654 4997 3688
rect 5031 3654 5043 3688
tri 5225 3669 5237 3681 se
rect 5237 3675 6292 3681
rect 5237 3669 5238 3675
rect 4317 3648 5043 3654
tri 5204 3648 5225 3669 se
rect 5225 3648 5238 3669
tri 5191 3635 5204 3648 se
rect 5204 3635 5238 3648
tri 5153 3597 5191 3635 se
rect 5191 3623 5238 3635
rect 5290 3623 5322 3675
rect 5374 3623 5406 3675
rect 5458 3669 6292 3675
rect 5458 3635 5675 3669
rect 5709 3635 6027 3669
rect 6061 3635 6292 3669
rect 5458 3623 6292 3635
rect 5191 3599 6292 3623
rect 5191 3597 5238 3599
tri 5119 3563 5153 3597 se
rect 5153 3563 5238 3597
tri 5109 3553 5119 3563 se
rect 5119 3553 5238 3563
rect -8872 3542 -8635 3548
rect -8872 3490 -8687 3542
rect -8872 3476 -8635 3490
rect -8872 3424 -8687 3476
rect -8872 3418 -8635 3424
rect 4057 3547 5238 3553
rect 5290 3547 5322 3599
rect 5374 3547 5406 3599
rect 5458 3597 6292 3599
rect 5458 3563 5675 3597
rect 5709 3563 6027 3597
rect 6061 3563 6292 3597
rect 5458 3547 6292 3563
rect 4057 3540 6292 3547
rect 4057 3506 4117 3540
rect 4151 3506 4821 3540
rect 4855 3523 6292 3540
rect 4855 3512 5238 3523
rect 5290 3512 5322 3523
rect 5374 3512 5406 3523
rect 5458 3512 6292 3523
rect 4855 3506 5126 3512
rect 4057 3478 5126 3506
rect 5160 3478 5198 3512
rect 5232 3478 5238 3512
rect 5304 3478 5322 3512
rect 5376 3478 5406 3512
rect 5458 3478 5486 3512
rect 5520 3478 5558 3512
rect 5592 3478 5630 3512
rect 5664 3478 5702 3512
rect 5736 3478 5774 3512
rect 5808 3478 5846 3512
rect 5880 3478 5918 3512
rect 5952 3478 5990 3512
rect 6024 3478 6062 3512
rect 6096 3478 6134 3512
rect 6168 3478 6206 3512
rect 6240 3478 6292 3512
rect 4057 3471 5238 3478
rect 5290 3471 5322 3478
rect 5374 3471 5406 3478
rect 5458 3471 6292 3478
rect 4057 3468 6292 3471
rect 4057 3434 4117 3468
rect 4151 3434 4821 3468
rect 4855 3448 6292 3468
rect 4855 3434 5238 3448
rect 4057 3396 5238 3434
rect 5290 3396 5322 3448
rect 5374 3396 5406 3448
rect 5458 3396 6292 3448
rect 4057 3390 6292 3396
tri -8913 3102 -8856 3159 se
rect -8856 3102 -8473 3159
rect -9284 2963 -8491 2964
rect -9329 2957 -8491 2963
rect -9329 2880 -8429 2957
rect -9329 2846 -8920 2880
rect -8886 2846 -8568 2880
rect -8534 2848 -8429 2880
tri -8429 2848 -8320 2957 nw
rect 4430 2899 4741 3074
rect -8534 2846 -8491 2848
rect -9329 2808 -8491 2846
rect -9329 2774 -8920 2808
rect -8886 2774 -8568 2808
rect -8534 2774 -8491 2808
tri -8491 2786 -8429 2848 nw
rect 6040 2842 6168 2848
rect 6092 2790 6116 2842
rect -9329 2761 -8491 2774
rect 6040 2776 6168 2790
rect 6092 2724 6116 2776
rect 6040 2718 6168 2724
rect -8750 2539 -8635 2545
rect -8750 2533 -8687 2539
rect -8750 2499 -8744 2533
rect -8710 2499 -8687 2533
rect -9012 2487 -8966 2499
rect -9012 2453 -9006 2487
rect -8972 2453 -8966 2487
rect -9012 2415 -8966 2453
rect -9012 2381 -9006 2415
rect -8972 2381 -8966 2415
rect -9012 2369 -8966 2381
rect -8833 2487 -8787 2499
rect -8833 2453 -8827 2487
rect -8793 2453 -8787 2487
rect -8833 2415 -8787 2453
rect -8750 2487 -8687 2499
rect 4316 2518 4387 2555
rect 5657 2525 5698 2569
rect 6220 2490 6294 2525
rect -8750 2473 -8635 2487
rect -8750 2461 -8687 2473
rect -8750 2427 -8744 2461
rect -8710 2427 -8687 2461
rect -8750 2421 -8687 2427
rect -8750 2415 -8635 2421
rect -8833 2381 -8827 2415
rect -8793 2381 -8787 2415
rect -8833 2369 -8787 2381
rect -9186 2343 -9140 2355
rect -9186 2309 -9180 2343
rect -9146 2309 -9140 2343
rect -9186 2271 -9140 2309
rect -9186 2237 -9180 2271
rect -9146 2237 -9140 2271
rect -9186 2225 -9140 2237
rect -9102 2336 -9056 2348
rect -9102 2302 -9096 2336
rect -9062 2302 -9056 2336
rect -8655 2336 -8609 2348
tri -9056 2302 -9052 2306 sw
rect -8655 2302 -8649 2336
rect -8615 2302 -8609 2336
rect -9102 2300 -9052 2302
tri -9052 2300 -9050 2302 sw
rect -9102 2264 -9050 2300
tri -9050 2264 -9014 2300 sw
tri -8691 2264 -8655 2300 se
rect -8655 2264 -8609 2302
rect -9102 2230 -9096 2264
rect -9062 2230 -8649 2264
rect -8615 2230 -8609 2264
rect -9102 2218 -8609 2230
rect 4310 2196 4377 2240
rect -9284 2129 -8491 2141
rect -9284 2095 -9272 2129
rect -9238 2095 -8920 2129
rect -8886 2095 -8491 2129
rect -9284 2079 -8491 2095
tri -8491 2079 -8429 2141 sw
rect -9284 2057 -8429 2079
rect -9284 2023 -9272 2057
rect -9238 2023 -8920 2057
rect -8886 2023 -8429 2057
rect -9284 2010 -8429 2023
tri -8429 2010 -8360 2079 sw
rect 5343 2073 5459 2079
rect -9284 1926 -8491 2010
rect 4346 1898 4513 2054
rect 5395 2021 5407 2073
rect 5343 2006 5459 2021
rect 5395 1954 5407 2006
rect 5343 1940 5459 1954
rect 5395 1888 5407 1940
rect 5343 1882 5459 1888
tri 6162 1847 6196 1881 ne
rect 6196 1744 6248 1881
tri 6248 1855 6274 1881 nw
rect 6003 1703 6045 1741
rect 6033 1340 6168 1457
<< via1 >>
rect 5099 7616 5151 7623
rect 5099 7582 5107 7616
rect 5107 7582 5141 7616
rect 5141 7582 5151 7616
rect 5099 7571 5151 7582
rect 5178 7616 5230 7623
rect 5256 7616 5308 7623
rect 5178 7582 5179 7616
rect 5179 7582 5213 7616
rect 5213 7582 5230 7616
rect 5256 7582 5285 7616
rect 5285 7582 5308 7616
rect 5178 7571 5230 7582
rect 5256 7571 5308 7582
rect 5099 7492 5151 7544
rect 5178 7492 5230 7544
rect 5256 7492 5308 7544
rect 5099 7413 5151 7465
rect 5178 7413 5230 7465
rect 5256 7413 5308 7465
rect 4434 7305 4486 7312
rect 4434 7271 4443 7305
rect 4443 7271 4477 7305
rect 4477 7271 4486 7305
rect 4434 7260 4486 7271
rect 4434 7233 4486 7245
rect 4434 7199 4443 7233
rect 4443 7199 4477 7233
rect 4477 7199 4486 7233
rect 4434 7193 4486 7199
rect 4603 7305 4655 7312
rect 4603 7271 4612 7305
rect 4612 7271 4646 7305
rect 4646 7271 4655 7305
rect 4603 7260 4655 7271
rect 4603 7233 4655 7245
rect 4603 7199 4612 7233
rect 4612 7199 4646 7233
rect 4646 7199 4655 7233
rect 4603 7193 4655 7199
rect 4786 7309 4838 7316
rect 4786 7275 4795 7309
rect 4795 7275 4829 7309
rect 4829 7275 4838 7309
rect 4786 7264 4838 7275
rect 4786 7237 4838 7249
rect 4786 7203 4795 7237
rect 4795 7203 4829 7237
rect 4829 7203 4838 7237
rect 4786 7197 4838 7203
rect 4959 7309 5011 7316
rect 4959 7275 4968 7309
rect 4968 7275 5002 7309
rect 5002 7275 5011 7309
rect 4959 7264 5011 7275
rect 4959 7237 5011 7249
rect 4959 7203 4968 7237
rect 4968 7203 5002 7237
rect 5002 7203 5011 7237
rect 4959 7197 5011 7203
rect 5436 7309 5488 7316
rect 5436 7275 5445 7309
rect 5445 7275 5479 7309
rect 5479 7275 5488 7309
rect 5436 7264 5488 7275
rect 5436 7237 5488 7249
rect 5436 7203 5445 7237
rect 5445 7203 5479 7237
rect 5479 7203 5488 7237
rect 5436 7197 5488 7203
rect 5659 7246 5711 7298
rect 5723 7246 5775 7298
rect 5442 7043 5494 7095
rect 5506 7043 5558 7095
rect 5002 6906 5054 6958
rect 5002 6842 5054 6894
rect 4695 6278 4747 6330
rect 4695 6214 4747 6266
rect 4786 6188 4838 6240
rect 4786 6124 4838 6176
rect 5002 6221 5054 6227
rect 5002 6187 5007 6221
rect 5007 6187 5041 6221
rect 5041 6187 5054 6221
rect 5002 6175 5054 6187
rect 5002 6149 5054 6161
rect 5002 6115 5007 6149
rect 5007 6115 5041 6149
rect 5041 6115 5054 6149
rect 5002 6109 5054 6115
rect 4821 6024 4873 6076
rect 4885 6024 4937 6076
rect 5729 6022 5781 6033
rect 4519 5939 4571 5991
rect 4519 5873 4571 5925
rect 5356 5924 5408 5976
rect 5356 5860 5408 5912
rect 5520 5941 5572 5993
rect 5520 5877 5572 5929
rect 5729 5988 5737 6022
rect 5737 5988 5771 6022
rect 5771 5988 5781 6022
rect 5729 5981 5781 5988
rect 5729 5950 5781 5962
rect 5729 5916 5737 5950
rect 5737 5916 5771 5950
rect 5771 5916 5781 5950
rect 5729 5910 5781 5916
rect 5095 5767 5147 5819
rect 5178 5811 5230 5819
rect 5178 5777 5183 5811
rect 5183 5777 5217 5811
rect 5217 5777 5230 5811
rect 5178 5767 5230 5777
rect 5261 5767 5313 5819
rect 5095 5701 5147 5753
rect 5178 5739 5230 5753
rect 5178 5705 5183 5739
rect 5183 5705 5217 5739
rect 5217 5705 5230 5739
rect 5178 5701 5230 5705
rect 5261 5701 5313 5753
rect 5095 5654 5147 5687
rect 5178 5654 5230 5687
rect 5261 5654 5313 5687
rect 5095 5635 5104 5654
rect 5104 5635 5138 5654
rect 5138 5635 5147 5654
rect 5178 5635 5210 5654
rect 5210 5635 5230 5654
rect 5261 5635 5282 5654
rect 5282 5635 5313 5654
rect 5095 5620 5104 5621
rect 5104 5620 5138 5621
rect 5138 5620 5147 5621
rect 5178 5620 5210 5621
rect 5210 5620 5230 5621
rect 5261 5620 5282 5621
rect 5282 5620 5313 5621
rect 5095 5569 5147 5620
rect 5178 5569 5230 5620
rect 5261 5569 5313 5620
rect 5095 5503 5147 5555
rect 5178 5503 5230 5555
rect 5261 5503 5313 5555
rect 5095 5437 5147 5489
rect 5178 5437 5230 5489
rect 5261 5437 5313 5489
rect 5095 5372 5147 5424
rect 5178 5372 5230 5424
rect 5261 5372 5313 5424
rect 3822 5271 3874 5323
rect 3886 5271 3938 5323
rect 4434 5046 4486 5098
rect 4434 4982 4486 5034
rect 4534 4937 4586 4989
rect 4598 4937 4650 4989
rect 5436 5045 5488 5051
rect 5436 5011 5469 5045
rect 5469 5011 5488 5045
rect 5436 4999 5488 5011
rect 5436 4973 5488 4985
rect 5436 4939 5469 4973
rect 5469 4939 5488 4973
rect 5436 4933 5488 4939
rect 5520 4860 5572 4912
rect 4565 4796 4617 4848
rect 4629 4796 4681 4848
rect 5520 4796 5572 4848
rect 5733 4788 5785 4840
rect 5733 4722 5785 4774
rect 6109 4246 6161 4252
rect 6109 4212 6116 4246
rect 6116 4212 6150 4246
rect 6150 4212 6161 4246
rect 6109 4200 6161 4212
rect 6109 4174 6161 4183
rect 6109 4140 6116 4174
rect 6116 4140 6150 4174
rect 6150 4140 6161 4174
rect 6109 4131 6161 4140
rect 3952 3910 4004 3962
rect 3952 3846 4004 3898
rect 4364 3829 4416 3881
rect 4428 3829 4480 3881
rect 4891 3824 4943 3876
rect 4891 3760 4943 3812
rect 5814 3885 5866 3891
rect 5814 3851 5850 3885
rect 5850 3851 5866 3885
rect 5814 3839 5866 3851
rect 5814 3813 5866 3825
rect 5814 3779 5850 3813
rect 5850 3779 5866 3813
rect 5814 3773 5866 3779
rect 5238 3623 5290 3675
rect 5322 3669 5374 3675
rect 5322 3635 5323 3669
rect 5323 3635 5357 3669
rect 5357 3635 5374 3669
rect 5322 3623 5374 3635
rect 5406 3623 5458 3675
rect -8687 3490 -8635 3542
rect -8687 3424 -8635 3476
rect 5238 3547 5290 3599
rect 5322 3597 5374 3599
rect 5322 3563 5323 3597
rect 5323 3563 5357 3597
rect 5357 3563 5374 3597
rect 5322 3547 5374 3563
rect 5406 3547 5458 3599
rect 5238 3512 5290 3523
rect 5322 3512 5374 3523
rect 5406 3512 5458 3523
rect 5238 3478 5270 3512
rect 5270 3478 5290 3512
rect 5322 3478 5342 3512
rect 5342 3478 5374 3512
rect 5406 3478 5414 3512
rect 5414 3478 5448 3512
rect 5448 3478 5458 3512
rect 5238 3471 5290 3478
rect 5322 3471 5374 3478
rect 5406 3471 5458 3478
rect 5238 3396 5290 3448
rect 5322 3396 5374 3448
rect 5406 3396 5458 3448
rect 6040 2790 6092 2842
rect 6116 2790 6168 2842
rect 6040 2724 6092 2776
rect 6116 2724 6168 2776
rect -8687 2487 -8635 2539
rect -8687 2421 -8635 2473
rect 5343 2021 5395 2073
rect 5407 2021 5459 2073
rect 5343 1954 5395 2006
rect 5407 1954 5459 2006
rect 5343 1888 5395 1940
rect 5407 1888 5459 1940
<< metal2 >>
rect 5093 7623 5314 7624
rect 5093 7571 5099 7623
rect 5151 7571 5178 7623
rect 5230 7571 5256 7623
rect 5308 7571 5314 7623
rect 5093 7544 5314 7571
rect 5093 7492 5099 7544
rect 5151 7492 5178 7544
rect 5230 7492 5256 7544
rect 5308 7492 5314 7544
tri 3907 5372 3952 5417 se
rect 3952 5372 4004 7362
tri 3858 5323 3907 5372 se
rect 3907 5323 4004 5372
rect 3816 5271 3822 5323
rect 3874 5271 3886 5323
rect 3938 5271 4004 5323
tri 3858 5177 3952 5271 ne
rect 3952 3962 4004 5271
rect 4434 7312 4486 7432
rect 4434 7245 4486 7260
rect 4434 5098 4486 7193
rect 4519 5991 4571 7453
rect 4519 5925 4571 5939
rect 4519 5867 4571 5873
rect 4603 7312 4655 7425
rect 4603 7245 4655 7260
tri 4590 5051 4603 5064 se
rect 4603 5051 4655 7193
rect 4786 7316 4838 7473
rect 4786 7249 4838 7264
rect 4959 7316 5011 7473
rect 4959 7249 5011 7264
tri 4925 7209 4959 7243 se
rect 4434 5034 4486 5046
tri 4538 4999 4590 5051 se
rect 4590 4999 4655 5051
rect 3952 3898 4004 3910
tri 4385 3891 4434 3940 se
rect 4434 3891 4486 4982
tri 4528 4989 4538 4999 se
rect 4538 4989 4655 4999
rect 4695 6330 4747 6336
rect 4695 6266 4747 6278
tri 4655 4989 4656 4990 sw
rect 4528 4937 4534 4989
rect 4586 4937 4598 4989
rect 4650 4937 4656 4989
tri 4655 4860 4695 4900 se
rect 4695 4860 4747 6214
rect 4786 6240 4838 7197
rect 4786 6176 4838 6188
rect 4786 6118 4838 6124
rect 4891 7197 4959 7209
rect 4891 7157 5011 7197
rect 5093 7465 5314 7492
rect 5093 7413 5099 7465
rect 5151 7413 5178 7465
rect 5230 7413 5256 7465
rect 5308 7413 5314 7465
tri 4890 6109 4891 6110 se
rect 4891 6109 4943 7157
tri 4943 7123 4977 7157 nw
tri 4857 6076 4890 6109 se
rect 4890 6076 4943 6109
rect 5002 6958 5054 6964
rect 5002 6894 5054 6906
rect 5002 6227 5054 6842
rect 5002 6161 5054 6175
rect 5002 6103 5054 6109
rect 4815 6024 4821 6076
rect 4873 6024 4885 6076
rect 4937 6024 4943 6076
tri 4857 5993 4888 6024 ne
rect 4888 5993 4943 6024
tri 4888 5990 4891 5993 ne
tri 4643 4848 4655 4860 se
rect 4655 4848 4747 4860
rect 4559 4796 4565 4848
rect 4617 4796 4629 4848
rect 4681 4796 4747 4848
tri 4376 3882 4385 3891 se
rect 4385 3882 4486 3891
tri 4375 3881 4376 3882 se
rect 4376 3881 4486 3882
rect 3952 3840 4004 3846
rect 4358 3829 4364 3881
rect 4416 3829 4428 3881
rect 4480 3829 4486 3881
rect 4891 3876 4943 5993
rect 4891 3812 4943 3824
rect 4891 3754 4943 3760
rect 5093 5819 5314 7413
rect 5436 7316 5488 7473
tri 5414 7264 5436 7286 se
tri 5399 7249 5414 7264 se
rect 5414 7249 5488 7264
tri 5380 7230 5399 7249 se
rect 5399 7230 5436 7249
rect 5356 7197 5436 7230
rect 5653 7246 5659 7298
rect 5711 7246 5723 7298
rect 5775 7246 5781 7298
tri 5695 7212 5729 7246 ne
rect 5356 7191 5488 7197
rect 5356 7157 5443 7191
tri 5443 7157 5477 7191 nw
rect 5356 7123 5409 7157
tri 5409 7123 5443 7157 nw
rect 5356 5976 5408 7123
tri 5408 7122 5409 7123 nw
rect 5356 5912 5408 5924
rect 5356 5854 5408 5860
rect 5436 7043 5442 7095
rect 5494 7043 5506 7095
rect 5558 7043 5564 7095
rect 5093 5767 5095 5819
rect 5147 5767 5178 5819
rect 5230 5767 5261 5819
rect 5313 5767 5314 5819
rect 5093 5753 5314 5767
rect 5093 5701 5095 5753
rect 5147 5701 5178 5753
rect 5230 5701 5261 5753
rect 5313 5701 5314 5753
rect 5093 5687 5314 5701
rect 5093 5635 5095 5687
rect 5147 5635 5178 5687
rect 5230 5635 5261 5687
rect 5313 5635 5314 5687
rect 5093 5621 5314 5635
rect 5093 5569 5095 5621
rect 5147 5569 5178 5621
rect 5230 5569 5261 5621
rect 5313 5569 5314 5621
rect 5093 5555 5314 5569
rect 5093 5503 5095 5555
rect 5147 5503 5178 5555
rect 5230 5503 5261 5555
rect 5313 5503 5314 5555
rect 5093 5489 5314 5503
rect 5093 5437 5095 5489
rect 5147 5437 5178 5489
rect 5230 5437 5261 5489
rect 5313 5437 5314 5489
rect 5093 5424 5314 5437
rect 5093 5372 5095 5424
rect 5147 5372 5178 5424
rect 5230 5372 5261 5424
rect 5313 5372 5314 5424
rect 5093 3897 5314 5372
rect 5436 5051 5488 7043
tri 5488 7009 5522 7043 nw
rect 5729 6033 5781 7246
rect 5436 4985 5488 4999
rect 5436 4927 5488 4933
rect 5520 5993 5572 5999
rect 5520 5929 5572 5941
rect 5729 5962 5781 5981
rect 5729 5904 5781 5910
rect 5520 4912 5572 5877
rect 5520 4848 5572 4860
rect 5520 4790 5572 4796
rect 5733 4840 5785 4846
rect 5733 4774 5785 4788
rect 5733 4716 5785 4722
rect 6109 4252 6161 4258
rect 6109 4183 6161 4200
rect 6109 4125 6161 4131
tri 5314 3897 5399 3982 sw
rect 5093 3891 5399 3897
tri 5399 3891 5405 3897 sw
rect 5814 3891 5866 3897
rect 5093 3839 5405 3891
tri 5405 3839 5457 3891 sw
rect 5093 3837 5457 3839
tri 5457 3837 5459 3839 sw
rect 5093 3675 5459 3837
rect 5814 3825 5866 3839
rect 5814 3767 5866 3773
rect 5093 3623 5238 3675
rect 5290 3623 5322 3675
rect 5374 3623 5406 3675
rect 5458 3623 5459 3675
rect 5093 3599 5459 3623
rect -8687 3542 -8635 3548
rect -8687 3476 -8635 3490
rect -8687 2539 -8635 3424
rect 5093 3547 5238 3599
rect 5290 3547 5322 3599
rect 5374 3547 5406 3599
rect 5458 3547 5459 3599
rect 5093 3523 5459 3547
rect 5093 3471 5238 3523
rect 5290 3471 5322 3523
rect 5374 3471 5406 3523
rect 5458 3471 5459 3523
rect 5093 3448 5459 3471
rect 5093 3396 5238 3448
rect 5290 3396 5322 3448
rect 5374 3396 5406 3448
rect 5458 3396 5459 3448
rect 5093 3310 5459 3396
tri 5093 3201 5202 3310 ne
rect 5202 3107 5459 3310
rect -8687 2473 -8635 2487
rect -8687 2415 -8635 2421
rect 5237 2073 5459 3107
rect 6040 2842 6168 2848
rect 6092 2790 6116 2842
rect 6040 2776 6168 2790
rect 6092 2724 6116 2776
rect 6040 2688 6168 2724
tri 5755 2254 5789 2288 se
rect 5237 2021 5343 2073
rect 5395 2021 5407 2073
rect 5237 2006 5459 2021
rect 5237 1954 5343 2006
rect 5395 1954 5407 2006
rect 5237 1940 5459 1954
rect 5237 1888 5343 1940
rect 5395 1888 5407 1940
rect 5237 1878 5459 1888
use sky130_fd_io__com_ctl_ls_octl  sky130_fd_io__com_ctl_ls_octl_0
timestamp 1688980957
transform 1 0 4281 0 -1 3202
box -71 10 2077 2019
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1688980957
transform -1 0 5943 0 1 5584
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1688980957
transform 1 0 5926 0 -1 5526
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_2
timestamp 1688980957
transform -1 0 5943 0 -1 7652
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_3
timestamp 1688980957
transform 1 0 5274 0 -1 5526
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_4
timestamp 1688980957
transform 1 0 5953 0 1 3442
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_0
timestamp 1688980957
transform -1 0 6295 0 1 5584
box 107 226 460 873
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_1
timestamp 1688980957
transform 1 0 5761 0 -1 7652
box 107 226 460 873
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_2
timestamp 1688980957
transform 1 0 5601 0 1 3442
box 107 226 460 873
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_3
timestamp 1688980957
transform 1 0 5574 0 -1 5526
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1688980957
transform 1 0 -8994 0 1 1902
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1688980957
transform -1 0 5291 0 1 5584
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_2
timestamp 1688980957
transform 1 0 5109 0 1 5584
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_3
timestamp 1688980957
transform 1 0 4281 0 1 5584
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_4
timestamp 1688980957
transform -1 0 4339 0 -1 7652
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_5
timestamp 1688980957
transform 1 0 4633 0 -1 7652
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_6
timestamp 1688980957
transform -1 0 5643 0 -1 7652
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_7
timestamp 1688980957
transform -1 0 4815 0 -1 7652
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1688980957
transform -1 0 -8812 0 1 1902
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1688980957
transform -1 0 4339 0 1 5584
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_2
timestamp 1688980957
transform -1 0 5783 0 1 3442
box 107 226 460 873
use sky130_fd_io__hvsbt_xor  sky130_fd_io__hvsbt_xor_0
timestamp 1688980957
transform 1 0 3805 0 -1 5656
box 213 167 1215 838
use sky130_fd_io__hvsbt_xorv2  sky130_fd_io__hvsbt_xorv2_0
timestamp 1688980957
transform 1 0 3772 0 1 3247
box 213 167 1215 838
<< labels >>
flabel metal2 s 4436 7368 4485 7431 3 FreeSans 520 270 0 0 DM_H[0]
port 2 nsew
flabel metal2 s 3965 7295 3991 7344 3 FreeSans 520 270 0 0 DM_H[2]
port 3 nsew
flabel metal2 s 5442 7419 5486 7468 3 FreeSans 520 270 0 0 DM_H_N[0]
port 4 nsew
flabel metal2 s 4968 7412 5002 7461 3 FreeSans 520 270 0 0 DM_H_N[1]
port 5 nsew
flabel metal2 s 4796 7417 4831 7462 3 FreeSans 520 270 0 0 DM_H_N[2]
port 6 nsew
flabel metal2 s 5020 6773 5051 6867 3 FreeSans 520 0 0 0 PUEN_2OR1_H
port 7 nsew
flabel metal2 s 4604 7370 4653 7423 3 FreeSans 520 270 0 0 DM_H[1]
port 1 nsew
flabel comment s 5456 7513 5456 7513 0 FreeSans 440 90 0 0 DM_H_N<0>
flabel comment s 4980 7575 4980 7575 0 FreeSans 440 270 0 0 DM_H_N<1>
flabel comment s 4804 7579 4804 7579 0 FreeSans 440 270 0 0 DM_H_N<2>
flabel comment s 4452 6892 4452 6892 0 FreeSans 440 90 0 0 DM_H<0>
flabel comment s 4630 6909 4630 6909 0 FreeSans 440 90 0 0 DM_H<1>
flabel comment s 3971 6510 3971 6510 0 FreeSans 440 270 0 0 DM_H<2>
flabel metal1 s 6014 6884 6044 6944 3 FreeSans 520 0 0 0 PDEN_H_N[1]
port 8 nsew
flabel metal1 s 6012 6289 6046 6353 3 FreeSans 520 0 0 0 PDEN_H_N[0]
port 9 nsew
flabel metal1 s 6003 1703 6045 1741 3 FreeSans 520 180 0 0 OD_H
port 10 nsew
flabel metal1 s 6220 2490 6294 2525 3 FreeSans 520 180 0 0 SLOW
port 11 nsew
flabel metal1 s 4316 2518 4387 2555 3 FreeSans 520 180 0 0 SLOW_H
port 12 nsew
flabel metal1 s 4310 2196 4377 2240 3 FreeSans 520 180 0 0 SLOW_H_N
port 13 nsew
flabel metal1 s 5657 2525 5698 2569 3 FreeSans 520 180 0 0 HLD_I_H_N
port 14 nsew
flabel metal1 s 5876 6498 6187 6730 3 FreeSans 520 0 0 0 VCC_IO
port 16 nsew
flabel metal1 s 6019 7436 6186 7606 3 FreeSans 520 0 0 0 VGND
port 15 nsew
flabel metal1 s 6033 1340 6168 1457 3 FreeSans 520 180 0 0 VPWR
port 17 nsew
flabel metal1 s 5876 4387 6187 4619 3 FreeSans 520 0 0 0 VCC_IO
port 16 nsew
flabel metal1 s 6019 5485 6186 5641 3 FreeSans 520 0 0 0 VGND
port 15 nsew
flabel metal1 s 6046 3453 6213 3609 3 FreeSans 520 0 0 0 VGND
port 15 nsew
flabel metal1 s 4346 1898 4513 2054 3 FreeSans 520 180 0 0 VGND
port 15 nsew
flabel metal1 s 4430 2899 4741 3074 3 FreeSans 520 180 0 0 VCC_IO
port 16 nsew
<< properties >>
string GDS_END 6893798
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6828852
<< end >>
