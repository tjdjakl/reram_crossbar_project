magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 439 203
rect 30 -17 64 21
<< locali >>
rect 103 333 169 493
rect 271 333 337 493
rect 103 299 443 333
rect 17 215 169 265
rect 203 215 353 265
rect 387 181 443 299
rect 271 131 443 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 17 299 69 527
rect 203 367 237 527
rect 371 367 422 527
rect 17 143 237 177
rect 17 51 85 143
rect 119 17 153 109
rect 187 93 237 143
rect 355 93 421 97
rect 187 51 421 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 203 215 353 265 6 A
port 1 nsew signal input
rlabel locali s 17 215 169 265 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 439 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 271 131 443 181 6 Y
port 7 nsew signal output
rlabel locali s 387 181 443 299 6 Y
port 7 nsew signal output
rlabel locali s 103 299 443 333 6 Y
port 7 nsew signal output
rlabel locali s 271 333 337 493 6 Y
port 7 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1636318
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1631338
<< end >>
