magic
tech sky130B
magscale 1 2
timestamp 1688980957
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1688980957
transform -1 0 16 0 1 13
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1688980957
transform 1 0 284 0 1 13
box 0 0 1 1
<< properties >>
string GDS_END 3728824
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3728342
<< end >>
