magic
tech sky130B
timestamp 1700618825
<< locali >>
rect 7895 3602 7954 8099
rect 6566 3515 9283 3602
rect 7895 -982 7954 3515
<< metal1 >>
rect 7895 7053 7960 7190
rect 7899 6034 7960 7053
rect 7895 5897 7960 6034
rect 7899 4895 7960 5897
rect 7895 4758 7960 4895
rect 6855 2469 6916 3762
rect 7204 2469 7265 3762
rect 7551 2469 7612 3762
rect 7899 3739 7960 4758
rect 7895 3602 7960 3739
rect 7899 2606 7960 3602
rect 7895 2469 7960 2606
rect 8243 2469 8304 3762
rect 8592 2469 8653 3762
rect 8939 2469 9000 3762
rect 7899 1450 7960 2469
rect 7895 1313 7960 1450
rect 7899 311 7960 1313
rect 7895 174 7960 311
rect 7899 -845 7960 174
rect 6580 -972 6680 -872
rect 7895 -982 7960 -845
<< metal2 >>
rect 6510 7237 6610 7337
rect 7534 7251 7957 7323
rect 6510 6081 6610 6181
rect 7534 6096 7957 6168
rect 6510 4942 6610 5042
rect 7533 4956 7956 5028
rect 6510 3786 6610 3886
rect 7529 3801 7952 3873
rect 6510 2653 6610 2753
rect 7531 2667 7954 2739
rect 6510 1497 6610 1597
rect 7531 1512 7954 1584
rect 6510 358 6610 458
rect 7527 372 7950 444
rect 6510 -798 6610 -698
rect 7539 -783 7962 -711
<< metal3 >>
rect 6599 8082 6699 8182
rect 6732 8082 6832 8182
rect 6946 8082 7046 8182
rect 7079 8082 7179 8182
rect 7295 8082 7395 8182
rect 7428 8082 7528 8182
rect 7642 8082 7742 8182
rect 7775 8082 7875 8182
rect 7987 8082 8087 8182
rect 8120 8082 8220 8182
rect 8334 8082 8434 8182
rect 8467 8082 8567 8182
rect 8683 8082 8783 8182
rect 8816 8082 8916 8182
rect 9030 8082 9130 8182
rect 9163 8082 9263 8182
rect 6608 3542 6687 4741
rect 6740 97 6820 8082
rect 6955 3541 7034 4740
rect 7087 96 7167 8082
rect 7304 3544 7383 4743
rect 7436 96 7516 8082
rect 7651 3544 7730 4743
rect 7783 97 7863 8082
rect 7996 3548 8075 4747
rect 8128 96 8208 8082
rect 8343 3542 8422 4741
rect 8475 96 8555 8082
rect 8692 3543 8771 4742
rect 8824 97 8904 8082
rect 9039 3544 9118 4743
rect 9171 96 9251 8082
use 16T16R  x1
timestamp 1700618825
transform 1 0 5821 0 1 3302
box 689 300 2074 4880
use 16T16R  x2
timestamp 1700618825
transform 1 0 5821 0 1 -1282
box 689 300 2074 4880
use 16T16R  x3
timestamp 1700618825
transform 1 0 7209 0 1 -1282
box 689 300 2074 4880
use 16T16R  x4
timestamp 1700618825
transform 1 0 7209 0 1 3302
box 689 300 2074 4880
<< labels >>
flabel metal3 9030 8082 9130 8182 0 FreeSans 128 0 0 0 SL8
port 25 nsew
flabel metal3 8683 8082 8783 8182 0 FreeSans 128 0 0 0 SL7
port 24 nsew
flabel metal3 8334 8082 8434 8182 0 FreeSans 128 0 0 0 SL6
port 23 nsew
flabel metal3 7987 8082 8087 8182 0 FreeSans 128 0 0 0 SL5
port 22 nsew
flabel metal3 7642 8082 7742 8182 0 FreeSans 128 0 0 0 SL4
port 20 nsew
flabel metal3 6946 8082 7046 8182 0 FreeSans 128 0 0 0 SL2
port 18 nsew
flabel metal3 6599 8082 6699 8182 0 FreeSans 128 0 0 0 SL1
port 17 nsew
flabel metal2 6510 -798 6610 -698 0 FreeSans 128 0 0 0 WL8
port 8 nsew
flabel metal2 6510 358 6610 458 0 FreeSans 128 0 0 0 WL7
port 7 nsew
flabel metal2 6510 1497 6610 1597 0 FreeSans 128 0 0 0 WL6
port 6 nsew
flabel metal2 6510 2653 6610 2753 0 FreeSans 128 0 0 0 WL5
port 5 nsew
flabel metal2 6510 3786 6610 3886 0 FreeSans 128 0 0 0 WL4
port 4 nsew
flabel metal2 6510 4942 6610 5042 0 FreeSans 128 0 0 0 WL3
port 3 nsew
flabel metal2 6510 6081 6610 6181 0 FreeSans 128 0 0 0 WL2
port 2 nsew
flabel metal2 6510 7237 6610 7337 0 FreeSans 128 0 0 0 WL1
port 1 nsew
flabel metal1 6580 -972 6680 -872 0 FreeSans 128 0 0 0 VSS
port 0 nsew
rlabel metal3 7295 8082 7395 8182 1 SL3
port 26 n
flabel metal3 9163 8082 9263 8182 0 FreeSans 128 0 0 0 BL8
port 16 nsew
flabel metal3 8816 8082 8916 8182 0 FreeSans 128 0 0 0 BL7
port 15 nsew
flabel metal3 8467 8082 8567 8182 0 FreeSans 128 0 0 0 BL6
port 14 nsew
flabel metal3 8120 8082 8220 8182 0 FreeSans 128 0 0 0 BL5
port 13 nsew
flabel metal3 7775 8082 7875 8182 0 FreeSans 128 0 0 0 BL4
port 12 nsew
flabel metal3 7428 8082 7528 8182 0 FreeSans 128 0 0 0 BL3
port 11 nsew
flabel metal3 7079 8082 7179 8182 0 FreeSans 128 0 0 0 BL2
port 10 nsew
flabel metal3 6732 8082 6832 8182 0 FreeSans 128 0 0 0 BL1
port 9 nsew
<< end >>
