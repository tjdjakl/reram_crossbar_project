magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect -38 261 222 582
<< pwell >>
rect 5 13 183 203
rect 29 -17 63 13
<< locali >>
rect 17 51 167 493
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 184 561
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 184 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 29 -17 63 17
rect 121 -17 155 17
<< metal1 >>
rect 0 561 184 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 184 561
rect 0 496 184 527
rect 0 17 184 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 184 17
rect 0 -48 184 -17
<< labels >>
rlabel locali s 17 51 167 493 6 DIODE
port 1 nsew signal input
rlabel metal1 s 0 -48 184 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 13 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 5 13 183 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 222 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 184 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 184 544
string LEFclass CORE ANTENNACELL
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2637356
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2633926
<< end >>
