magic
tech sky130B
magscale 1 2
timestamp 1700618825
<< pwell >>
rect -1225 -2133 1225 2133
<< psubdiff >>
rect -1189 2063 -1093 2097
rect 1093 2063 1189 2097
rect -1189 2001 -1155 2063
rect 1155 2001 1189 2063
rect -1189 -2063 -1155 -2001
rect 1155 -2063 1189 -2001
rect -1189 -2097 -1093 -2063
rect 1093 -2097 1189 -2063
<< psubdiffcont >>
rect -1093 2063 1093 2097
rect -1189 -2001 -1155 2001
rect 1155 -2001 1189 2001
rect -1093 -2097 1093 -2063
<< poly >>
rect -1059 -1917 -993 -1537
rect -1059 -1951 -1043 -1917
rect -1009 -1951 -993 -1917
rect -1059 -1967 -993 -1951
rect 993 -1917 1059 -1537
rect 993 -1951 1009 -1917
rect 1043 -1951 1059 -1917
rect 993 -1967 1059 -1951
<< polycont >>
rect -1043 -1951 -1009 -1917
rect 1009 -1951 1043 -1917
<< npolyres >>
rect -1059 1901 -885 1967
rect -1059 -1537 -993 1901
rect -951 -1367 -885 1901
rect -843 1901 -669 1967
rect -843 -1367 -777 1901
rect -951 -1433 -777 -1367
rect -735 -1367 -669 1901
rect -627 1901 -453 1967
rect -627 -1367 -561 1901
rect -735 -1433 -561 -1367
rect -519 -1367 -453 1901
rect -411 1901 -237 1967
rect -411 -1367 -345 1901
rect -519 -1433 -345 -1367
rect -303 -1367 -237 1901
rect -195 1901 -21 1967
rect -195 -1367 -129 1901
rect -303 -1433 -129 -1367
rect -87 -1367 -21 1901
rect 21 1901 195 1967
rect 21 -1367 87 1901
rect -87 -1433 87 -1367
rect 129 -1367 195 1901
rect 237 1901 411 1967
rect 237 -1367 303 1901
rect 129 -1433 303 -1367
rect 345 -1367 411 1901
rect 453 1901 627 1967
rect 453 -1367 519 1901
rect 345 -1433 519 -1367
rect 561 -1367 627 1901
rect 669 1901 843 1967
rect 669 -1367 735 1901
rect 561 -1433 735 -1367
rect 777 -1367 843 1901
rect 885 1901 1059 1967
rect 885 -1367 951 1901
rect 777 -1433 951 -1367
rect 993 -1537 1059 1901
<< locali >>
rect -1189 2063 -1093 2097
rect 1093 2063 1189 2097
rect -1189 2001 -1155 2063
rect 1155 2001 1189 2063
rect -1059 -1951 -1043 -1917
rect -1009 -1951 -993 -1917
rect 993 -1951 1009 -1917
rect 1043 -1951 1059 -1917
rect -1189 -2063 -1155 -2001
rect 1155 -2063 1189 -2001
rect -1189 -2097 -1093 -2063
rect 1093 -2097 1189 -2063
<< properties >>
string FIXED_BBOX -1172 -2080 1172 2080
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.330 l 17 m 1 nx 20 wmin 0.330 lmin 1.650 rho 48.2 val 51.686k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 1 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
