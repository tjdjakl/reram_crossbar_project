magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< pwell >>
rect 15 163 2283 1225
<< mvnmos >>
rect 241 189 341 1199
rect 397 189 497 1199
rect 553 189 653 1199
rect 709 189 809 1199
rect 865 189 965 1199
rect 1021 189 1121 1199
rect 1177 189 1277 1199
rect 1333 189 1433 1199
rect 1489 189 1589 1199
rect 1645 189 1745 1199
rect 1801 189 1901 1199
rect 1957 189 2057 1199
<< mvndiff >>
rect 181 1187 241 1199
rect 181 1153 196 1187
rect 230 1153 241 1187
rect 181 1119 241 1153
rect 181 1085 196 1119
rect 230 1085 241 1119
rect 181 1051 241 1085
rect 181 1017 196 1051
rect 230 1017 241 1051
rect 181 983 241 1017
rect 181 949 196 983
rect 230 949 241 983
rect 181 915 241 949
rect 181 881 196 915
rect 230 881 241 915
rect 181 847 241 881
rect 181 813 196 847
rect 230 813 241 847
rect 181 779 241 813
rect 181 745 196 779
rect 230 745 241 779
rect 181 711 241 745
rect 181 677 196 711
rect 230 677 241 711
rect 181 643 241 677
rect 181 609 196 643
rect 230 609 241 643
rect 181 575 241 609
rect 181 541 196 575
rect 230 541 241 575
rect 181 507 241 541
rect 181 473 196 507
rect 230 473 241 507
rect 181 439 241 473
rect 181 405 196 439
rect 230 405 241 439
rect 181 371 241 405
rect 181 337 196 371
rect 230 337 241 371
rect 181 303 241 337
rect 181 269 196 303
rect 230 269 241 303
rect 181 235 241 269
rect 181 201 196 235
rect 230 201 241 235
rect 181 189 241 201
rect 341 1187 397 1199
rect 341 1153 352 1187
rect 386 1153 397 1187
rect 341 1119 397 1153
rect 341 1085 352 1119
rect 386 1085 397 1119
rect 341 1051 397 1085
rect 341 1017 352 1051
rect 386 1017 397 1051
rect 341 983 397 1017
rect 341 949 352 983
rect 386 949 397 983
rect 341 915 397 949
rect 341 881 352 915
rect 386 881 397 915
rect 341 847 397 881
rect 341 813 352 847
rect 386 813 397 847
rect 341 779 397 813
rect 341 745 352 779
rect 386 745 397 779
rect 341 711 397 745
rect 341 677 352 711
rect 386 677 397 711
rect 341 643 397 677
rect 341 609 352 643
rect 386 609 397 643
rect 341 575 397 609
rect 341 541 352 575
rect 386 541 397 575
rect 341 507 397 541
rect 341 473 352 507
rect 386 473 397 507
rect 341 439 397 473
rect 341 405 352 439
rect 386 405 397 439
rect 341 371 397 405
rect 341 337 352 371
rect 386 337 397 371
rect 341 303 397 337
rect 341 269 352 303
rect 386 269 397 303
rect 341 235 397 269
rect 341 201 352 235
rect 386 201 397 235
rect 341 189 397 201
rect 497 1187 553 1199
rect 497 1153 508 1187
rect 542 1153 553 1187
rect 497 1119 553 1153
rect 497 1085 508 1119
rect 542 1085 553 1119
rect 497 1051 553 1085
rect 497 1017 508 1051
rect 542 1017 553 1051
rect 497 983 553 1017
rect 497 949 508 983
rect 542 949 553 983
rect 497 915 553 949
rect 497 881 508 915
rect 542 881 553 915
rect 497 847 553 881
rect 497 813 508 847
rect 542 813 553 847
rect 497 779 553 813
rect 497 745 508 779
rect 542 745 553 779
rect 497 711 553 745
rect 497 677 508 711
rect 542 677 553 711
rect 497 643 553 677
rect 497 609 508 643
rect 542 609 553 643
rect 497 575 553 609
rect 497 541 508 575
rect 542 541 553 575
rect 497 507 553 541
rect 497 473 508 507
rect 542 473 553 507
rect 497 439 553 473
rect 497 405 508 439
rect 542 405 553 439
rect 497 371 553 405
rect 497 337 508 371
rect 542 337 553 371
rect 497 303 553 337
rect 497 269 508 303
rect 542 269 553 303
rect 497 235 553 269
rect 497 201 508 235
rect 542 201 553 235
rect 497 189 553 201
rect 653 1187 709 1199
rect 653 1153 664 1187
rect 698 1153 709 1187
rect 653 1119 709 1153
rect 653 1085 664 1119
rect 698 1085 709 1119
rect 653 1051 709 1085
rect 653 1017 664 1051
rect 698 1017 709 1051
rect 653 983 709 1017
rect 653 949 664 983
rect 698 949 709 983
rect 653 915 709 949
rect 653 881 664 915
rect 698 881 709 915
rect 653 847 709 881
rect 653 813 664 847
rect 698 813 709 847
rect 653 779 709 813
rect 653 745 664 779
rect 698 745 709 779
rect 653 711 709 745
rect 653 677 664 711
rect 698 677 709 711
rect 653 643 709 677
rect 653 609 664 643
rect 698 609 709 643
rect 653 575 709 609
rect 653 541 664 575
rect 698 541 709 575
rect 653 507 709 541
rect 653 473 664 507
rect 698 473 709 507
rect 653 439 709 473
rect 653 405 664 439
rect 698 405 709 439
rect 653 371 709 405
rect 653 337 664 371
rect 698 337 709 371
rect 653 303 709 337
rect 653 269 664 303
rect 698 269 709 303
rect 653 235 709 269
rect 653 201 664 235
rect 698 201 709 235
rect 653 189 709 201
rect 809 1187 865 1199
rect 809 1153 820 1187
rect 854 1153 865 1187
rect 809 1119 865 1153
rect 809 1085 820 1119
rect 854 1085 865 1119
rect 809 1051 865 1085
rect 809 1017 820 1051
rect 854 1017 865 1051
rect 809 983 865 1017
rect 809 949 820 983
rect 854 949 865 983
rect 809 915 865 949
rect 809 881 820 915
rect 854 881 865 915
rect 809 847 865 881
rect 809 813 820 847
rect 854 813 865 847
rect 809 779 865 813
rect 809 745 820 779
rect 854 745 865 779
rect 809 711 865 745
rect 809 677 820 711
rect 854 677 865 711
rect 809 643 865 677
rect 809 609 820 643
rect 854 609 865 643
rect 809 575 865 609
rect 809 541 820 575
rect 854 541 865 575
rect 809 507 865 541
rect 809 473 820 507
rect 854 473 865 507
rect 809 439 865 473
rect 809 405 820 439
rect 854 405 865 439
rect 809 371 865 405
rect 809 337 820 371
rect 854 337 865 371
rect 809 303 865 337
rect 809 269 820 303
rect 854 269 865 303
rect 809 235 865 269
rect 809 201 820 235
rect 854 201 865 235
rect 809 189 865 201
rect 965 1187 1021 1199
rect 965 1153 976 1187
rect 1010 1153 1021 1187
rect 965 1119 1021 1153
rect 965 1085 976 1119
rect 1010 1085 1021 1119
rect 965 1051 1021 1085
rect 965 1017 976 1051
rect 1010 1017 1021 1051
rect 965 983 1021 1017
rect 965 949 976 983
rect 1010 949 1021 983
rect 965 915 1021 949
rect 965 881 976 915
rect 1010 881 1021 915
rect 965 847 1021 881
rect 965 813 976 847
rect 1010 813 1021 847
rect 965 779 1021 813
rect 965 745 976 779
rect 1010 745 1021 779
rect 965 711 1021 745
rect 965 677 976 711
rect 1010 677 1021 711
rect 965 643 1021 677
rect 965 609 976 643
rect 1010 609 1021 643
rect 965 575 1021 609
rect 965 541 976 575
rect 1010 541 1021 575
rect 965 507 1021 541
rect 965 473 976 507
rect 1010 473 1021 507
rect 965 439 1021 473
rect 965 405 976 439
rect 1010 405 1021 439
rect 965 371 1021 405
rect 965 337 976 371
rect 1010 337 1021 371
rect 965 303 1021 337
rect 965 269 976 303
rect 1010 269 1021 303
rect 965 235 1021 269
rect 965 201 976 235
rect 1010 201 1021 235
rect 965 189 1021 201
rect 1121 1187 1177 1199
rect 1121 1153 1132 1187
rect 1166 1153 1177 1187
rect 1121 1119 1177 1153
rect 1121 1085 1132 1119
rect 1166 1085 1177 1119
rect 1121 1051 1177 1085
rect 1121 1017 1132 1051
rect 1166 1017 1177 1051
rect 1121 983 1177 1017
rect 1121 949 1132 983
rect 1166 949 1177 983
rect 1121 915 1177 949
rect 1121 881 1132 915
rect 1166 881 1177 915
rect 1121 847 1177 881
rect 1121 813 1132 847
rect 1166 813 1177 847
rect 1121 779 1177 813
rect 1121 745 1132 779
rect 1166 745 1177 779
rect 1121 711 1177 745
rect 1121 677 1132 711
rect 1166 677 1177 711
rect 1121 643 1177 677
rect 1121 609 1132 643
rect 1166 609 1177 643
rect 1121 575 1177 609
rect 1121 541 1132 575
rect 1166 541 1177 575
rect 1121 507 1177 541
rect 1121 473 1132 507
rect 1166 473 1177 507
rect 1121 439 1177 473
rect 1121 405 1132 439
rect 1166 405 1177 439
rect 1121 371 1177 405
rect 1121 337 1132 371
rect 1166 337 1177 371
rect 1121 303 1177 337
rect 1121 269 1132 303
rect 1166 269 1177 303
rect 1121 235 1177 269
rect 1121 201 1132 235
rect 1166 201 1177 235
rect 1121 189 1177 201
rect 1277 1187 1333 1199
rect 1277 1153 1288 1187
rect 1322 1153 1333 1187
rect 1277 1119 1333 1153
rect 1277 1085 1288 1119
rect 1322 1085 1333 1119
rect 1277 1051 1333 1085
rect 1277 1017 1288 1051
rect 1322 1017 1333 1051
rect 1277 983 1333 1017
rect 1277 949 1288 983
rect 1322 949 1333 983
rect 1277 915 1333 949
rect 1277 881 1288 915
rect 1322 881 1333 915
rect 1277 847 1333 881
rect 1277 813 1288 847
rect 1322 813 1333 847
rect 1277 779 1333 813
rect 1277 745 1288 779
rect 1322 745 1333 779
rect 1277 711 1333 745
rect 1277 677 1288 711
rect 1322 677 1333 711
rect 1277 643 1333 677
rect 1277 609 1288 643
rect 1322 609 1333 643
rect 1277 575 1333 609
rect 1277 541 1288 575
rect 1322 541 1333 575
rect 1277 507 1333 541
rect 1277 473 1288 507
rect 1322 473 1333 507
rect 1277 439 1333 473
rect 1277 405 1288 439
rect 1322 405 1333 439
rect 1277 371 1333 405
rect 1277 337 1288 371
rect 1322 337 1333 371
rect 1277 303 1333 337
rect 1277 269 1288 303
rect 1322 269 1333 303
rect 1277 235 1333 269
rect 1277 201 1288 235
rect 1322 201 1333 235
rect 1277 189 1333 201
rect 1433 1187 1489 1199
rect 1433 1153 1444 1187
rect 1478 1153 1489 1187
rect 1433 1119 1489 1153
rect 1433 1085 1444 1119
rect 1478 1085 1489 1119
rect 1433 1051 1489 1085
rect 1433 1017 1444 1051
rect 1478 1017 1489 1051
rect 1433 983 1489 1017
rect 1433 949 1444 983
rect 1478 949 1489 983
rect 1433 915 1489 949
rect 1433 881 1444 915
rect 1478 881 1489 915
rect 1433 847 1489 881
rect 1433 813 1444 847
rect 1478 813 1489 847
rect 1433 779 1489 813
rect 1433 745 1444 779
rect 1478 745 1489 779
rect 1433 711 1489 745
rect 1433 677 1444 711
rect 1478 677 1489 711
rect 1433 643 1489 677
rect 1433 609 1444 643
rect 1478 609 1489 643
rect 1433 575 1489 609
rect 1433 541 1444 575
rect 1478 541 1489 575
rect 1433 507 1489 541
rect 1433 473 1444 507
rect 1478 473 1489 507
rect 1433 439 1489 473
rect 1433 405 1444 439
rect 1478 405 1489 439
rect 1433 371 1489 405
rect 1433 337 1444 371
rect 1478 337 1489 371
rect 1433 303 1489 337
rect 1433 269 1444 303
rect 1478 269 1489 303
rect 1433 235 1489 269
rect 1433 201 1444 235
rect 1478 201 1489 235
rect 1433 189 1489 201
rect 1589 1187 1645 1199
rect 1589 1153 1600 1187
rect 1634 1153 1645 1187
rect 1589 1119 1645 1153
rect 1589 1085 1600 1119
rect 1634 1085 1645 1119
rect 1589 1051 1645 1085
rect 1589 1017 1600 1051
rect 1634 1017 1645 1051
rect 1589 983 1645 1017
rect 1589 949 1600 983
rect 1634 949 1645 983
rect 1589 915 1645 949
rect 1589 881 1600 915
rect 1634 881 1645 915
rect 1589 847 1645 881
rect 1589 813 1600 847
rect 1634 813 1645 847
rect 1589 779 1645 813
rect 1589 745 1600 779
rect 1634 745 1645 779
rect 1589 711 1645 745
rect 1589 677 1600 711
rect 1634 677 1645 711
rect 1589 643 1645 677
rect 1589 609 1600 643
rect 1634 609 1645 643
rect 1589 575 1645 609
rect 1589 541 1600 575
rect 1634 541 1645 575
rect 1589 507 1645 541
rect 1589 473 1600 507
rect 1634 473 1645 507
rect 1589 439 1645 473
rect 1589 405 1600 439
rect 1634 405 1645 439
rect 1589 371 1645 405
rect 1589 337 1600 371
rect 1634 337 1645 371
rect 1589 303 1645 337
rect 1589 269 1600 303
rect 1634 269 1645 303
rect 1589 235 1645 269
rect 1589 201 1600 235
rect 1634 201 1645 235
rect 1589 189 1645 201
rect 1745 1187 1801 1199
rect 1745 1153 1756 1187
rect 1790 1153 1801 1187
rect 1745 1119 1801 1153
rect 1745 1085 1756 1119
rect 1790 1085 1801 1119
rect 1745 1051 1801 1085
rect 1745 1017 1756 1051
rect 1790 1017 1801 1051
rect 1745 983 1801 1017
rect 1745 949 1756 983
rect 1790 949 1801 983
rect 1745 915 1801 949
rect 1745 881 1756 915
rect 1790 881 1801 915
rect 1745 847 1801 881
rect 1745 813 1756 847
rect 1790 813 1801 847
rect 1745 779 1801 813
rect 1745 745 1756 779
rect 1790 745 1801 779
rect 1745 711 1801 745
rect 1745 677 1756 711
rect 1790 677 1801 711
rect 1745 643 1801 677
rect 1745 609 1756 643
rect 1790 609 1801 643
rect 1745 575 1801 609
rect 1745 541 1756 575
rect 1790 541 1801 575
rect 1745 507 1801 541
rect 1745 473 1756 507
rect 1790 473 1801 507
rect 1745 439 1801 473
rect 1745 405 1756 439
rect 1790 405 1801 439
rect 1745 371 1801 405
rect 1745 337 1756 371
rect 1790 337 1801 371
rect 1745 303 1801 337
rect 1745 269 1756 303
rect 1790 269 1801 303
rect 1745 235 1801 269
rect 1745 201 1756 235
rect 1790 201 1801 235
rect 1745 189 1801 201
rect 1901 1187 1957 1199
rect 1901 1153 1912 1187
rect 1946 1153 1957 1187
rect 1901 1119 1957 1153
rect 1901 1085 1912 1119
rect 1946 1085 1957 1119
rect 1901 1051 1957 1085
rect 1901 1017 1912 1051
rect 1946 1017 1957 1051
rect 1901 983 1957 1017
rect 1901 949 1912 983
rect 1946 949 1957 983
rect 1901 915 1957 949
rect 1901 881 1912 915
rect 1946 881 1957 915
rect 1901 847 1957 881
rect 1901 813 1912 847
rect 1946 813 1957 847
rect 1901 779 1957 813
rect 1901 745 1912 779
rect 1946 745 1957 779
rect 1901 711 1957 745
rect 1901 677 1912 711
rect 1946 677 1957 711
rect 1901 643 1957 677
rect 1901 609 1912 643
rect 1946 609 1957 643
rect 1901 575 1957 609
rect 1901 541 1912 575
rect 1946 541 1957 575
rect 1901 507 1957 541
rect 1901 473 1912 507
rect 1946 473 1957 507
rect 1901 439 1957 473
rect 1901 405 1912 439
rect 1946 405 1957 439
rect 1901 371 1957 405
rect 1901 337 1912 371
rect 1946 337 1957 371
rect 1901 303 1957 337
rect 1901 269 1912 303
rect 1946 269 1957 303
rect 1901 235 1957 269
rect 1901 201 1912 235
rect 1946 201 1957 235
rect 1901 189 1957 201
rect 2057 1187 2117 1199
rect 2057 1153 2068 1187
rect 2102 1153 2117 1187
rect 2057 1119 2117 1153
rect 2057 1085 2068 1119
rect 2102 1085 2117 1119
rect 2057 1051 2117 1085
rect 2057 1017 2068 1051
rect 2102 1017 2117 1051
rect 2057 983 2117 1017
rect 2057 949 2068 983
rect 2102 949 2117 983
rect 2057 915 2117 949
rect 2057 881 2068 915
rect 2102 881 2117 915
rect 2057 847 2117 881
rect 2057 813 2068 847
rect 2102 813 2117 847
rect 2057 779 2117 813
rect 2057 745 2068 779
rect 2102 745 2117 779
rect 2057 711 2117 745
rect 2057 677 2068 711
rect 2102 677 2117 711
rect 2057 643 2117 677
rect 2057 609 2068 643
rect 2102 609 2117 643
rect 2057 575 2117 609
rect 2057 541 2068 575
rect 2102 541 2117 575
rect 2057 507 2117 541
rect 2057 473 2068 507
rect 2102 473 2117 507
rect 2057 439 2117 473
rect 2057 405 2068 439
rect 2102 405 2117 439
rect 2057 371 2117 405
rect 2057 337 2068 371
rect 2102 337 2117 371
rect 2057 303 2117 337
rect 2057 269 2068 303
rect 2102 269 2117 303
rect 2057 235 2117 269
rect 2057 201 2068 235
rect 2102 201 2117 235
rect 2057 189 2117 201
<< mvndiffc >>
rect 196 1153 230 1187
rect 196 1085 230 1119
rect 196 1017 230 1051
rect 196 949 230 983
rect 196 881 230 915
rect 196 813 230 847
rect 196 745 230 779
rect 196 677 230 711
rect 196 609 230 643
rect 196 541 230 575
rect 196 473 230 507
rect 196 405 230 439
rect 196 337 230 371
rect 196 269 230 303
rect 196 201 230 235
rect 352 1153 386 1187
rect 352 1085 386 1119
rect 352 1017 386 1051
rect 352 949 386 983
rect 352 881 386 915
rect 352 813 386 847
rect 352 745 386 779
rect 352 677 386 711
rect 352 609 386 643
rect 352 541 386 575
rect 352 473 386 507
rect 352 405 386 439
rect 352 337 386 371
rect 352 269 386 303
rect 352 201 386 235
rect 508 1153 542 1187
rect 508 1085 542 1119
rect 508 1017 542 1051
rect 508 949 542 983
rect 508 881 542 915
rect 508 813 542 847
rect 508 745 542 779
rect 508 677 542 711
rect 508 609 542 643
rect 508 541 542 575
rect 508 473 542 507
rect 508 405 542 439
rect 508 337 542 371
rect 508 269 542 303
rect 508 201 542 235
rect 664 1153 698 1187
rect 664 1085 698 1119
rect 664 1017 698 1051
rect 664 949 698 983
rect 664 881 698 915
rect 664 813 698 847
rect 664 745 698 779
rect 664 677 698 711
rect 664 609 698 643
rect 664 541 698 575
rect 664 473 698 507
rect 664 405 698 439
rect 664 337 698 371
rect 664 269 698 303
rect 664 201 698 235
rect 820 1153 854 1187
rect 820 1085 854 1119
rect 820 1017 854 1051
rect 820 949 854 983
rect 820 881 854 915
rect 820 813 854 847
rect 820 745 854 779
rect 820 677 854 711
rect 820 609 854 643
rect 820 541 854 575
rect 820 473 854 507
rect 820 405 854 439
rect 820 337 854 371
rect 820 269 854 303
rect 820 201 854 235
rect 976 1153 1010 1187
rect 976 1085 1010 1119
rect 976 1017 1010 1051
rect 976 949 1010 983
rect 976 881 1010 915
rect 976 813 1010 847
rect 976 745 1010 779
rect 976 677 1010 711
rect 976 609 1010 643
rect 976 541 1010 575
rect 976 473 1010 507
rect 976 405 1010 439
rect 976 337 1010 371
rect 976 269 1010 303
rect 976 201 1010 235
rect 1132 1153 1166 1187
rect 1132 1085 1166 1119
rect 1132 1017 1166 1051
rect 1132 949 1166 983
rect 1132 881 1166 915
rect 1132 813 1166 847
rect 1132 745 1166 779
rect 1132 677 1166 711
rect 1132 609 1166 643
rect 1132 541 1166 575
rect 1132 473 1166 507
rect 1132 405 1166 439
rect 1132 337 1166 371
rect 1132 269 1166 303
rect 1132 201 1166 235
rect 1288 1153 1322 1187
rect 1288 1085 1322 1119
rect 1288 1017 1322 1051
rect 1288 949 1322 983
rect 1288 881 1322 915
rect 1288 813 1322 847
rect 1288 745 1322 779
rect 1288 677 1322 711
rect 1288 609 1322 643
rect 1288 541 1322 575
rect 1288 473 1322 507
rect 1288 405 1322 439
rect 1288 337 1322 371
rect 1288 269 1322 303
rect 1288 201 1322 235
rect 1444 1153 1478 1187
rect 1444 1085 1478 1119
rect 1444 1017 1478 1051
rect 1444 949 1478 983
rect 1444 881 1478 915
rect 1444 813 1478 847
rect 1444 745 1478 779
rect 1444 677 1478 711
rect 1444 609 1478 643
rect 1444 541 1478 575
rect 1444 473 1478 507
rect 1444 405 1478 439
rect 1444 337 1478 371
rect 1444 269 1478 303
rect 1444 201 1478 235
rect 1600 1153 1634 1187
rect 1600 1085 1634 1119
rect 1600 1017 1634 1051
rect 1600 949 1634 983
rect 1600 881 1634 915
rect 1600 813 1634 847
rect 1600 745 1634 779
rect 1600 677 1634 711
rect 1600 609 1634 643
rect 1600 541 1634 575
rect 1600 473 1634 507
rect 1600 405 1634 439
rect 1600 337 1634 371
rect 1600 269 1634 303
rect 1600 201 1634 235
rect 1756 1153 1790 1187
rect 1756 1085 1790 1119
rect 1756 1017 1790 1051
rect 1756 949 1790 983
rect 1756 881 1790 915
rect 1756 813 1790 847
rect 1756 745 1790 779
rect 1756 677 1790 711
rect 1756 609 1790 643
rect 1756 541 1790 575
rect 1756 473 1790 507
rect 1756 405 1790 439
rect 1756 337 1790 371
rect 1756 269 1790 303
rect 1756 201 1790 235
rect 1912 1153 1946 1187
rect 1912 1085 1946 1119
rect 1912 1017 1946 1051
rect 1912 949 1946 983
rect 1912 881 1946 915
rect 1912 813 1946 847
rect 1912 745 1946 779
rect 1912 677 1946 711
rect 1912 609 1946 643
rect 1912 541 1946 575
rect 1912 473 1946 507
rect 1912 405 1946 439
rect 1912 337 1946 371
rect 1912 269 1946 303
rect 1912 201 1946 235
rect 2068 1153 2102 1187
rect 2068 1085 2102 1119
rect 2068 1017 2102 1051
rect 2068 949 2102 983
rect 2068 881 2102 915
rect 2068 813 2102 847
rect 2068 745 2102 779
rect 2068 677 2102 711
rect 2068 609 2102 643
rect 2068 541 2102 575
rect 2068 473 2102 507
rect 2068 405 2102 439
rect 2068 337 2102 371
rect 2068 269 2102 303
rect 2068 201 2102 235
<< mvpsubdiff >>
rect 41 1187 181 1199
rect 41 201 60 1187
rect 162 201 181 1187
rect 41 189 181 201
rect 2117 1187 2257 1199
rect 2117 201 2136 1187
rect 2238 201 2257 1187
rect 2117 189 2257 201
<< mvpsubdiffcont >>
rect 60 201 162 1187
rect 2136 201 2238 1187
<< poly >>
rect 383 1367 1915 1388
rect 190 1275 341 1291
rect 190 1241 206 1275
rect 240 1241 341 1275
rect 383 1265 418 1367
rect 1880 1265 1915 1367
rect 383 1249 1915 1265
rect 1957 1275 2108 1291
rect 190 1225 341 1241
rect 241 1199 341 1225
rect 397 1199 497 1249
rect 553 1199 653 1249
rect 709 1199 809 1249
rect 865 1199 965 1249
rect 1021 1199 1121 1249
rect 1177 1199 1277 1249
rect 1333 1199 1433 1249
rect 1489 1199 1589 1249
rect 1645 1199 1745 1249
rect 1801 1199 1901 1249
rect 1957 1241 2058 1275
rect 2092 1241 2108 1275
rect 1957 1225 2108 1241
rect 1957 1199 2057 1225
rect 241 163 341 189
rect 190 147 341 163
rect 190 113 206 147
rect 240 113 341 147
rect 397 139 497 189
rect 553 139 653 189
rect 709 139 809 189
rect 865 139 965 189
rect 1021 139 1121 189
rect 1177 139 1277 189
rect 1333 139 1433 189
rect 1489 139 1589 189
rect 1645 139 1745 189
rect 1801 139 1901 189
rect 1957 163 2057 189
rect 1957 147 2108 163
rect 190 97 341 113
rect 383 123 1915 139
rect 383 21 418 123
rect 1880 21 1915 123
rect 1957 113 2058 147
rect 2092 113 2108 147
rect 1957 97 2108 113
rect 383 0 1915 21
<< polycont >>
rect 206 1241 240 1275
rect 418 1265 1880 1367
rect 2058 1241 2092 1275
rect 206 113 240 147
rect 418 21 1880 123
rect 2058 113 2092 147
<< locali >>
rect 385 1369 1913 1388
rect 190 1275 256 1291
rect 190 1241 206 1275
rect 240 1241 256 1275
rect 385 1263 412 1369
rect 1886 1263 1913 1369
rect 385 1251 1913 1263
rect 2042 1275 2108 1291
rect 190 1225 256 1241
rect 2042 1241 2058 1275
rect 2092 1241 2108 1275
rect 2042 1225 2108 1241
rect 190 1203 230 1225
rect 2068 1203 2108 1225
rect 41 1187 230 1203
rect 41 201 60 1187
rect 162 1153 196 1187
rect 162 1119 230 1153
rect 162 1085 196 1119
rect 162 1051 230 1085
rect 162 1017 196 1051
rect 162 983 230 1017
rect 162 949 196 983
rect 162 915 230 949
rect 162 881 196 915
rect 162 847 230 881
rect 162 813 196 847
rect 162 779 230 813
rect 162 745 196 779
rect 162 711 230 745
rect 162 677 196 711
rect 162 643 230 677
rect 162 609 196 643
rect 162 575 230 609
rect 162 541 196 575
rect 162 507 230 541
rect 162 473 196 507
rect 162 439 230 473
rect 162 405 196 439
rect 162 371 230 405
rect 162 337 196 371
rect 162 303 230 337
rect 162 269 196 303
rect 162 235 230 269
rect 162 201 196 235
rect 41 185 230 201
rect 352 1187 386 1203
rect 352 1119 386 1145
rect 352 1051 386 1073
rect 352 983 386 1001
rect 352 915 386 929
rect 352 847 386 857
rect 352 779 386 785
rect 352 711 386 713
rect 352 675 386 677
rect 352 603 386 609
rect 352 531 386 541
rect 352 459 386 473
rect 352 387 386 405
rect 352 315 386 337
rect 352 243 386 269
rect 352 185 386 201
rect 508 1187 542 1203
rect 508 1119 542 1145
rect 508 1051 542 1073
rect 508 983 542 1001
rect 508 915 542 929
rect 508 847 542 857
rect 508 779 542 785
rect 508 711 542 713
rect 508 675 542 677
rect 508 603 542 609
rect 508 531 542 541
rect 508 459 542 473
rect 508 387 542 405
rect 508 315 542 337
rect 508 243 542 269
rect 508 185 542 201
rect 664 1187 698 1203
rect 664 1119 698 1145
rect 664 1051 698 1073
rect 664 983 698 1001
rect 664 915 698 929
rect 664 847 698 857
rect 664 779 698 785
rect 664 711 698 713
rect 664 675 698 677
rect 664 603 698 609
rect 664 531 698 541
rect 664 459 698 473
rect 664 387 698 405
rect 664 315 698 337
rect 664 243 698 269
rect 664 185 698 201
rect 820 1187 854 1203
rect 820 1119 854 1145
rect 820 1051 854 1073
rect 820 983 854 1001
rect 820 915 854 929
rect 820 847 854 857
rect 820 779 854 785
rect 820 711 854 713
rect 820 675 854 677
rect 820 603 854 609
rect 820 531 854 541
rect 820 459 854 473
rect 820 387 854 405
rect 820 315 854 337
rect 820 243 854 269
rect 820 185 854 201
rect 976 1187 1010 1203
rect 976 1119 1010 1145
rect 976 1051 1010 1073
rect 976 983 1010 1001
rect 976 915 1010 929
rect 976 847 1010 857
rect 976 779 1010 785
rect 976 711 1010 713
rect 976 675 1010 677
rect 976 603 1010 609
rect 976 531 1010 541
rect 976 459 1010 473
rect 976 387 1010 405
rect 976 315 1010 337
rect 976 243 1010 269
rect 976 185 1010 201
rect 1132 1187 1166 1203
rect 1132 1119 1166 1145
rect 1132 1051 1166 1073
rect 1132 983 1166 1001
rect 1132 915 1166 929
rect 1132 847 1166 857
rect 1132 779 1166 785
rect 1132 711 1166 713
rect 1132 675 1166 677
rect 1132 603 1166 609
rect 1132 531 1166 541
rect 1132 459 1166 473
rect 1132 387 1166 405
rect 1132 315 1166 337
rect 1132 243 1166 269
rect 1132 185 1166 201
rect 1288 1187 1322 1203
rect 1288 1119 1322 1145
rect 1288 1051 1322 1073
rect 1288 983 1322 1001
rect 1288 915 1322 929
rect 1288 847 1322 857
rect 1288 779 1322 785
rect 1288 711 1322 713
rect 1288 675 1322 677
rect 1288 603 1322 609
rect 1288 531 1322 541
rect 1288 459 1322 473
rect 1288 387 1322 405
rect 1288 315 1322 337
rect 1288 243 1322 269
rect 1288 185 1322 201
rect 1444 1187 1478 1203
rect 1444 1119 1478 1145
rect 1444 1051 1478 1073
rect 1444 983 1478 1001
rect 1444 915 1478 929
rect 1444 847 1478 857
rect 1444 779 1478 785
rect 1444 711 1478 713
rect 1444 675 1478 677
rect 1444 603 1478 609
rect 1444 531 1478 541
rect 1444 459 1478 473
rect 1444 387 1478 405
rect 1444 315 1478 337
rect 1444 243 1478 269
rect 1444 185 1478 201
rect 1600 1187 1634 1203
rect 1600 1119 1634 1145
rect 1600 1051 1634 1073
rect 1600 983 1634 1001
rect 1600 915 1634 929
rect 1600 847 1634 857
rect 1600 779 1634 785
rect 1600 711 1634 713
rect 1600 675 1634 677
rect 1600 603 1634 609
rect 1600 531 1634 541
rect 1600 459 1634 473
rect 1600 387 1634 405
rect 1600 315 1634 337
rect 1600 243 1634 269
rect 1600 185 1634 201
rect 1756 1187 1790 1203
rect 1756 1119 1790 1145
rect 1756 1051 1790 1073
rect 1756 983 1790 1001
rect 1756 915 1790 929
rect 1756 847 1790 857
rect 1756 779 1790 785
rect 1756 711 1790 713
rect 1756 675 1790 677
rect 1756 603 1790 609
rect 1756 531 1790 541
rect 1756 459 1790 473
rect 1756 387 1790 405
rect 1756 315 1790 337
rect 1756 243 1790 269
rect 1756 185 1790 201
rect 1912 1187 1946 1203
rect 1912 1119 1946 1145
rect 1912 1051 1946 1073
rect 1912 983 1946 1001
rect 1912 915 1946 929
rect 1912 847 1946 857
rect 1912 779 1946 785
rect 1912 711 1946 713
rect 1912 675 1946 677
rect 1912 603 1946 609
rect 1912 531 1946 541
rect 1912 459 1946 473
rect 1912 387 1946 405
rect 1912 315 1946 337
rect 1912 243 1946 269
rect 1912 185 1946 201
rect 2068 1187 2257 1203
rect 2102 1153 2136 1187
rect 2068 1119 2136 1153
rect 2102 1085 2136 1119
rect 2068 1051 2136 1085
rect 2102 1017 2136 1051
rect 2068 983 2136 1017
rect 2102 949 2136 983
rect 2068 915 2136 949
rect 2102 881 2136 915
rect 2068 847 2136 881
rect 2102 813 2136 847
rect 2068 779 2136 813
rect 2102 745 2136 779
rect 2068 711 2136 745
rect 2102 677 2136 711
rect 2068 643 2136 677
rect 2102 609 2136 643
rect 2068 575 2136 609
rect 2102 541 2136 575
rect 2068 507 2136 541
rect 2102 473 2136 507
rect 2068 439 2136 473
rect 2102 405 2136 439
rect 2068 371 2136 405
rect 2102 337 2136 371
rect 2068 303 2136 337
rect 2102 269 2136 303
rect 2068 235 2136 269
rect 2102 201 2136 235
rect 2238 201 2257 1187
rect 2068 185 2257 201
rect 190 163 230 185
rect 2068 163 2108 185
rect 190 147 256 163
rect 190 113 206 147
rect 240 113 256 147
rect 2042 147 2108 163
rect 190 97 256 113
rect 385 125 1913 137
rect 385 19 412 125
rect 1886 19 1913 125
rect 2042 113 2058 147
rect 2092 113 2108 147
rect 2042 97 2108 113
rect 385 0 1913 19
<< viali >>
rect 412 1367 1886 1369
rect 412 1265 418 1367
rect 418 1265 1880 1367
rect 1880 1265 1886 1367
rect 412 1263 1886 1265
rect 60 1145 94 1179
rect 60 1073 94 1107
rect 60 1001 94 1035
rect 60 929 94 963
rect 60 857 94 891
rect 60 785 94 819
rect 60 713 94 747
rect 60 641 94 675
rect 60 569 94 603
rect 60 497 94 531
rect 60 425 94 459
rect 60 353 94 387
rect 60 281 94 315
rect 60 209 94 243
rect 352 1153 386 1179
rect 352 1145 386 1153
rect 352 1085 386 1107
rect 352 1073 386 1085
rect 352 1017 386 1035
rect 352 1001 386 1017
rect 352 949 386 963
rect 352 929 386 949
rect 352 881 386 891
rect 352 857 386 881
rect 352 813 386 819
rect 352 785 386 813
rect 352 745 386 747
rect 352 713 386 745
rect 352 643 386 675
rect 352 641 386 643
rect 352 575 386 603
rect 352 569 386 575
rect 352 507 386 531
rect 352 497 386 507
rect 352 439 386 459
rect 352 425 386 439
rect 352 371 386 387
rect 352 353 386 371
rect 352 303 386 315
rect 352 281 386 303
rect 352 235 386 243
rect 352 209 386 235
rect 508 1153 542 1179
rect 508 1145 542 1153
rect 508 1085 542 1107
rect 508 1073 542 1085
rect 508 1017 542 1035
rect 508 1001 542 1017
rect 508 949 542 963
rect 508 929 542 949
rect 508 881 542 891
rect 508 857 542 881
rect 508 813 542 819
rect 508 785 542 813
rect 508 745 542 747
rect 508 713 542 745
rect 508 643 542 675
rect 508 641 542 643
rect 508 575 542 603
rect 508 569 542 575
rect 508 507 542 531
rect 508 497 542 507
rect 508 439 542 459
rect 508 425 542 439
rect 508 371 542 387
rect 508 353 542 371
rect 508 303 542 315
rect 508 281 542 303
rect 508 235 542 243
rect 508 209 542 235
rect 664 1153 698 1179
rect 664 1145 698 1153
rect 664 1085 698 1107
rect 664 1073 698 1085
rect 664 1017 698 1035
rect 664 1001 698 1017
rect 664 949 698 963
rect 664 929 698 949
rect 664 881 698 891
rect 664 857 698 881
rect 664 813 698 819
rect 664 785 698 813
rect 664 745 698 747
rect 664 713 698 745
rect 664 643 698 675
rect 664 641 698 643
rect 664 575 698 603
rect 664 569 698 575
rect 664 507 698 531
rect 664 497 698 507
rect 664 439 698 459
rect 664 425 698 439
rect 664 371 698 387
rect 664 353 698 371
rect 664 303 698 315
rect 664 281 698 303
rect 664 235 698 243
rect 664 209 698 235
rect 820 1153 854 1179
rect 820 1145 854 1153
rect 820 1085 854 1107
rect 820 1073 854 1085
rect 820 1017 854 1035
rect 820 1001 854 1017
rect 820 949 854 963
rect 820 929 854 949
rect 820 881 854 891
rect 820 857 854 881
rect 820 813 854 819
rect 820 785 854 813
rect 820 745 854 747
rect 820 713 854 745
rect 820 643 854 675
rect 820 641 854 643
rect 820 575 854 603
rect 820 569 854 575
rect 820 507 854 531
rect 820 497 854 507
rect 820 439 854 459
rect 820 425 854 439
rect 820 371 854 387
rect 820 353 854 371
rect 820 303 854 315
rect 820 281 854 303
rect 820 235 854 243
rect 820 209 854 235
rect 976 1153 1010 1179
rect 976 1145 1010 1153
rect 976 1085 1010 1107
rect 976 1073 1010 1085
rect 976 1017 1010 1035
rect 976 1001 1010 1017
rect 976 949 1010 963
rect 976 929 1010 949
rect 976 881 1010 891
rect 976 857 1010 881
rect 976 813 1010 819
rect 976 785 1010 813
rect 976 745 1010 747
rect 976 713 1010 745
rect 976 643 1010 675
rect 976 641 1010 643
rect 976 575 1010 603
rect 976 569 1010 575
rect 976 507 1010 531
rect 976 497 1010 507
rect 976 439 1010 459
rect 976 425 1010 439
rect 976 371 1010 387
rect 976 353 1010 371
rect 976 303 1010 315
rect 976 281 1010 303
rect 976 235 1010 243
rect 976 209 1010 235
rect 1132 1153 1166 1179
rect 1132 1145 1166 1153
rect 1132 1085 1166 1107
rect 1132 1073 1166 1085
rect 1132 1017 1166 1035
rect 1132 1001 1166 1017
rect 1132 949 1166 963
rect 1132 929 1166 949
rect 1132 881 1166 891
rect 1132 857 1166 881
rect 1132 813 1166 819
rect 1132 785 1166 813
rect 1132 745 1166 747
rect 1132 713 1166 745
rect 1132 643 1166 675
rect 1132 641 1166 643
rect 1132 575 1166 603
rect 1132 569 1166 575
rect 1132 507 1166 531
rect 1132 497 1166 507
rect 1132 439 1166 459
rect 1132 425 1166 439
rect 1132 371 1166 387
rect 1132 353 1166 371
rect 1132 303 1166 315
rect 1132 281 1166 303
rect 1132 235 1166 243
rect 1132 209 1166 235
rect 1288 1153 1322 1179
rect 1288 1145 1322 1153
rect 1288 1085 1322 1107
rect 1288 1073 1322 1085
rect 1288 1017 1322 1035
rect 1288 1001 1322 1017
rect 1288 949 1322 963
rect 1288 929 1322 949
rect 1288 881 1322 891
rect 1288 857 1322 881
rect 1288 813 1322 819
rect 1288 785 1322 813
rect 1288 745 1322 747
rect 1288 713 1322 745
rect 1288 643 1322 675
rect 1288 641 1322 643
rect 1288 575 1322 603
rect 1288 569 1322 575
rect 1288 507 1322 531
rect 1288 497 1322 507
rect 1288 439 1322 459
rect 1288 425 1322 439
rect 1288 371 1322 387
rect 1288 353 1322 371
rect 1288 303 1322 315
rect 1288 281 1322 303
rect 1288 235 1322 243
rect 1288 209 1322 235
rect 1444 1153 1478 1179
rect 1444 1145 1478 1153
rect 1444 1085 1478 1107
rect 1444 1073 1478 1085
rect 1444 1017 1478 1035
rect 1444 1001 1478 1017
rect 1444 949 1478 963
rect 1444 929 1478 949
rect 1444 881 1478 891
rect 1444 857 1478 881
rect 1444 813 1478 819
rect 1444 785 1478 813
rect 1444 745 1478 747
rect 1444 713 1478 745
rect 1444 643 1478 675
rect 1444 641 1478 643
rect 1444 575 1478 603
rect 1444 569 1478 575
rect 1444 507 1478 531
rect 1444 497 1478 507
rect 1444 439 1478 459
rect 1444 425 1478 439
rect 1444 371 1478 387
rect 1444 353 1478 371
rect 1444 303 1478 315
rect 1444 281 1478 303
rect 1444 235 1478 243
rect 1444 209 1478 235
rect 1600 1153 1634 1179
rect 1600 1145 1634 1153
rect 1600 1085 1634 1107
rect 1600 1073 1634 1085
rect 1600 1017 1634 1035
rect 1600 1001 1634 1017
rect 1600 949 1634 963
rect 1600 929 1634 949
rect 1600 881 1634 891
rect 1600 857 1634 881
rect 1600 813 1634 819
rect 1600 785 1634 813
rect 1600 745 1634 747
rect 1600 713 1634 745
rect 1600 643 1634 675
rect 1600 641 1634 643
rect 1600 575 1634 603
rect 1600 569 1634 575
rect 1600 507 1634 531
rect 1600 497 1634 507
rect 1600 439 1634 459
rect 1600 425 1634 439
rect 1600 371 1634 387
rect 1600 353 1634 371
rect 1600 303 1634 315
rect 1600 281 1634 303
rect 1600 235 1634 243
rect 1600 209 1634 235
rect 1756 1153 1790 1179
rect 1756 1145 1790 1153
rect 1756 1085 1790 1107
rect 1756 1073 1790 1085
rect 1756 1017 1790 1035
rect 1756 1001 1790 1017
rect 1756 949 1790 963
rect 1756 929 1790 949
rect 1756 881 1790 891
rect 1756 857 1790 881
rect 1756 813 1790 819
rect 1756 785 1790 813
rect 1756 745 1790 747
rect 1756 713 1790 745
rect 1756 643 1790 675
rect 1756 641 1790 643
rect 1756 575 1790 603
rect 1756 569 1790 575
rect 1756 507 1790 531
rect 1756 497 1790 507
rect 1756 439 1790 459
rect 1756 425 1790 439
rect 1756 371 1790 387
rect 1756 353 1790 371
rect 1756 303 1790 315
rect 1756 281 1790 303
rect 1756 235 1790 243
rect 1756 209 1790 235
rect 1912 1153 1946 1179
rect 1912 1145 1946 1153
rect 1912 1085 1946 1107
rect 1912 1073 1946 1085
rect 1912 1017 1946 1035
rect 1912 1001 1946 1017
rect 1912 949 1946 963
rect 1912 929 1946 949
rect 1912 881 1946 891
rect 1912 857 1946 881
rect 1912 813 1946 819
rect 1912 785 1946 813
rect 1912 745 1946 747
rect 1912 713 1946 745
rect 1912 643 1946 675
rect 1912 641 1946 643
rect 1912 575 1946 603
rect 1912 569 1946 575
rect 1912 507 1946 531
rect 1912 497 1946 507
rect 1912 439 1946 459
rect 1912 425 1946 439
rect 1912 371 1946 387
rect 1912 353 1946 371
rect 1912 303 1946 315
rect 1912 281 1946 303
rect 1912 235 1946 243
rect 1912 209 1946 235
rect 2204 1145 2238 1179
rect 2204 1073 2238 1107
rect 2204 1001 2238 1035
rect 2204 929 2238 963
rect 2204 857 2238 891
rect 2204 785 2238 819
rect 2204 713 2238 747
rect 2204 641 2238 675
rect 2204 569 2238 603
rect 2204 497 2238 531
rect 2204 425 2238 459
rect 2204 353 2238 387
rect 2204 281 2238 315
rect 2204 209 2238 243
rect 412 123 1886 125
rect 412 21 418 123
rect 418 21 1880 123
rect 1880 21 1886 123
rect 412 19 1886 21
<< metal1 >>
rect 381 1369 1917 1388
rect 381 1263 412 1369
rect 1886 1263 1917 1369
rect 381 1251 1917 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 343 1179 395 1191
rect 343 1145 352 1179
rect 386 1145 395 1179
rect 343 1107 395 1145
rect 343 1073 352 1107
rect 386 1073 395 1107
rect 343 1035 395 1073
rect 343 1001 352 1035
rect 386 1001 395 1035
rect 343 963 395 1001
rect 343 929 352 963
rect 386 929 395 963
rect 343 891 395 929
rect 343 857 352 891
rect 386 857 395 891
rect 343 819 395 857
rect 343 785 352 819
rect 386 785 395 819
rect 343 747 395 785
rect 343 713 352 747
rect 386 713 395 747
rect 343 675 395 713
rect 343 641 352 675
rect 386 641 395 675
rect 343 639 395 641
rect 343 575 352 587
rect 386 575 395 587
rect 343 511 352 523
rect 386 511 395 523
rect 343 447 352 459
rect 386 447 395 459
rect 343 387 395 395
rect 343 383 352 387
rect 386 383 395 387
rect 343 319 395 331
rect 343 255 395 267
rect 343 197 395 203
rect 499 1185 551 1191
rect 499 1121 551 1133
rect 499 1057 551 1069
rect 499 1001 508 1005
rect 542 1001 551 1005
rect 499 993 551 1001
rect 499 929 508 941
rect 542 929 551 941
rect 499 865 508 877
rect 542 865 551 877
rect 499 801 508 813
rect 542 801 551 813
rect 499 747 551 749
rect 499 713 508 747
rect 542 713 551 747
rect 499 675 551 713
rect 499 641 508 675
rect 542 641 551 675
rect 499 603 551 641
rect 499 569 508 603
rect 542 569 551 603
rect 499 531 551 569
rect 499 497 508 531
rect 542 497 551 531
rect 499 459 551 497
rect 499 425 508 459
rect 542 425 551 459
rect 499 387 551 425
rect 499 353 508 387
rect 542 353 551 387
rect 499 315 551 353
rect 499 281 508 315
rect 542 281 551 315
rect 499 243 551 281
rect 499 209 508 243
rect 542 209 551 243
rect 499 197 551 209
rect 655 1179 707 1191
rect 655 1145 664 1179
rect 698 1145 707 1179
rect 655 1107 707 1145
rect 655 1073 664 1107
rect 698 1073 707 1107
rect 655 1035 707 1073
rect 655 1001 664 1035
rect 698 1001 707 1035
rect 655 963 707 1001
rect 655 929 664 963
rect 698 929 707 963
rect 655 891 707 929
rect 655 857 664 891
rect 698 857 707 891
rect 655 819 707 857
rect 655 785 664 819
rect 698 785 707 819
rect 655 747 707 785
rect 655 713 664 747
rect 698 713 707 747
rect 655 675 707 713
rect 655 641 664 675
rect 698 641 707 675
rect 655 639 707 641
rect 655 575 664 587
rect 698 575 707 587
rect 655 511 664 523
rect 698 511 707 523
rect 655 447 664 459
rect 698 447 707 459
rect 655 387 707 395
rect 655 383 664 387
rect 698 383 707 387
rect 655 319 707 331
rect 655 255 707 267
rect 655 197 707 203
rect 811 1185 863 1191
rect 811 1121 863 1133
rect 811 1057 863 1069
rect 811 1001 820 1005
rect 854 1001 863 1005
rect 811 993 863 1001
rect 811 929 820 941
rect 854 929 863 941
rect 811 865 820 877
rect 854 865 863 877
rect 811 801 820 813
rect 854 801 863 813
rect 811 747 863 749
rect 811 713 820 747
rect 854 713 863 747
rect 811 675 863 713
rect 811 641 820 675
rect 854 641 863 675
rect 811 603 863 641
rect 811 569 820 603
rect 854 569 863 603
rect 811 531 863 569
rect 811 497 820 531
rect 854 497 863 531
rect 811 459 863 497
rect 811 425 820 459
rect 854 425 863 459
rect 811 387 863 425
rect 811 353 820 387
rect 854 353 863 387
rect 811 315 863 353
rect 811 281 820 315
rect 854 281 863 315
rect 811 243 863 281
rect 811 209 820 243
rect 854 209 863 243
rect 811 197 863 209
rect 967 1179 1019 1191
rect 967 1145 976 1179
rect 1010 1145 1019 1179
rect 967 1107 1019 1145
rect 967 1073 976 1107
rect 1010 1073 1019 1107
rect 967 1035 1019 1073
rect 967 1001 976 1035
rect 1010 1001 1019 1035
rect 967 963 1019 1001
rect 967 929 976 963
rect 1010 929 1019 963
rect 967 891 1019 929
rect 967 857 976 891
rect 1010 857 1019 891
rect 967 819 1019 857
rect 967 785 976 819
rect 1010 785 1019 819
rect 967 747 1019 785
rect 967 713 976 747
rect 1010 713 1019 747
rect 967 675 1019 713
rect 967 641 976 675
rect 1010 641 1019 675
rect 967 639 1019 641
rect 967 575 976 587
rect 1010 575 1019 587
rect 967 511 976 523
rect 1010 511 1019 523
rect 967 447 976 459
rect 1010 447 1019 459
rect 967 387 1019 395
rect 967 383 976 387
rect 1010 383 1019 387
rect 967 319 1019 331
rect 967 255 1019 267
rect 967 197 1019 203
rect 1123 1185 1175 1191
rect 1123 1121 1175 1133
rect 1123 1057 1175 1069
rect 1123 1001 1132 1005
rect 1166 1001 1175 1005
rect 1123 993 1175 1001
rect 1123 929 1132 941
rect 1166 929 1175 941
rect 1123 865 1132 877
rect 1166 865 1175 877
rect 1123 801 1132 813
rect 1166 801 1175 813
rect 1123 747 1175 749
rect 1123 713 1132 747
rect 1166 713 1175 747
rect 1123 675 1175 713
rect 1123 641 1132 675
rect 1166 641 1175 675
rect 1123 603 1175 641
rect 1123 569 1132 603
rect 1166 569 1175 603
rect 1123 531 1175 569
rect 1123 497 1132 531
rect 1166 497 1175 531
rect 1123 459 1175 497
rect 1123 425 1132 459
rect 1166 425 1175 459
rect 1123 387 1175 425
rect 1123 353 1132 387
rect 1166 353 1175 387
rect 1123 315 1175 353
rect 1123 281 1132 315
rect 1166 281 1175 315
rect 1123 243 1175 281
rect 1123 209 1132 243
rect 1166 209 1175 243
rect 1123 197 1175 209
rect 1279 1179 1331 1191
rect 1279 1145 1288 1179
rect 1322 1145 1331 1179
rect 1279 1107 1331 1145
rect 1279 1073 1288 1107
rect 1322 1073 1331 1107
rect 1279 1035 1331 1073
rect 1279 1001 1288 1035
rect 1322 1001 1331 1035
rect 1279 963 1331 1001
rect 1279 929 1288 963
rect 1322 929 1331 963
rect 1279 891 1331 929
rect 1279 857 1288 891
rect 1322 857 1331 891
rect 1279 819 1331 857
rect 1279 785 1288 819
rect 1322 785 1331 819
rect 1279 747 1331 785
rect 1279 713 1288 747
rect 1322 713 1331 747
rect 1279 675 1331 713
rect 1279 641 1288 675
rect 1322 641 1331 675
rect 1279 639 1331 641
rect 1279 575 1288 587
rect 1322 575 1331 587
rect 1279 511 1288 523
rect 1322 511 1331 523
rect 1279 447 1288 459
rect 1322 447 1331 459
rect 1279 387 1331 395
rect 1279 383 1288 387
rect 1322 383 1331 387
rect 1279 319 1331 331
rect 1279 255 1331 267
rect 1279 197 1331 203
rect 1435 1185 1487 1191
rect 1435 1121 1487 1133
rect 1435 1057 1487 1069
rect 1435 1001 1444 1005
rect 1478 1001 1487 1005
rect 1435 993 1487 1001
rect 1435 929 1444 941
rect 1478 929 1487 941
rect 1435 865 1444 877
rect 1478 865 1487 877
rect 1435 801 1444 813
rect 1478 801 1487 813
rect 1435 747 1487 749
rect 1435 713 1444 747
rect 1478 713 1487 747
rect 1435 675 1487 713
rect 1435 641 1444 675
rect 1478 641 1487 675
rect 1435 603 1487 641
rect 1435 569 1444 603
rect 1478 569 1487 603
rect 1435 531 1487 569
rect 1435 497 1444 531
rect 1478 497 1487 531
rect 1435 459 1487 497
rect 1435 425 1444 459
rect 1478 425 1487 459
rect 1435 387 1487 425
rect 1435 353 1444 387
rect 1478 353 1487 387
rect 1435 315 1487 353
rect 1435 281 1444 315
rect 1478 281 1487 315
rect 1435 243 1487 281
rect 1435 209 1444 243
rect 1478 209 1487 243
rect 1435 197 1487 209
rect 1591 1179 1643 1191
rect 1591 1145 1600 1179
rect 1634 1145 1643 1179
rect 1591 1107 1643 1145
rect 1591 1073 1600 1107
rect 1634 1073 1643 1107
rect 1591 1035 1643 1073
rect 1591 1001 1600 1035
rect 1634 1001 1643 1035
rect 1591 963 1643 1001
rect 1591 929 1600 963
rect 1634 929 1643 963
rect 1591 891 1643 929
rect 1591 857 1600 891
rect 1634 857 1643 891
rect 1591 819 1643 857
rect 1591 785 1600 819
rect 1634 785 1643 819
rect 1591 747 1643 785
rect 1591 713 1600 747
rect 1634 713 1643 747
rect 1591 675 1643 713
rect 1591 641 1600 675
rect 1634 641 1643 675
rect 1591 639 1643 641
rect 1591 575 1600 587
rect 1634 575 1643 587
rect 1591 511 1600 523
rect 1634 511 1643 523
rect 1591 447 1600 459
rect 1634 447 1643 459
rect 1591 387 1643 395
rect 1591 383 1600 387
rect 1634 383 1643 387
rect 1591 319 1643 331
rect 1591 255 1643 267
rect 1591 197 1643 203
rect 1747 1185 1799 1191
rect 1747 1121 1799 1133
rect 1747 1057 1799 1069
rect 1747 1001 1756 1005
rect 1790 1001 1799 1005
rect 1747 993 1799 1001
rect 1747 929 1756 941
rect 1790 929 1799 941
rect 1747 865 1756 877
rect 1790 865 1799 877
rect 1747 801 1756 813
rect 1790 801 1799 813
rect 1747 747 1799 749
rect 1747 713 1756 747
rect 1790 713 1799 747
rect 1747 675 1799 713
rect 1747 641 1756 675
rect 1790 641 1799 675
rect 1747 603 1799 641
rect 1747 569 1756 603
rect 1790 569 1799 603
rect 1747 531 1799 569
rect 1747 497 1756 531
rect 1790 497 1799 531
rect 1747 459 1799 497
rect 1747 425 1756 459
rect 1790 425 1799 459
rect 1747 387 1799 425
rect 1747 353 1756 387
rect 1790 353 1799 387
rect 1747 315 1799 353
rect 1747 281 1756 315
rect 1790 281 1799 315
rect 1747 243 1799 281
rect 1747 209 1756 243
rect 1790 209 1799 243
rect 1747 197 1799 209
rect 1903 1179 1955 1191
rect 1903 1145 1912 1179
rect 1946 1145 1955 1179
rect 1903 1107 1955 1145
rect 1903 1073 1912 1107
rect 1946 1073 1955 1107
rect 1903 1035 1955 1073
rect 1903 1001 1912 1035
rect 1946 1001 1955 1035
rect 1903 963 1955 1001
rect 1903 929 1912 963
rect 1946 929 1955 963
rect 1903 891 1955 929
rect 1903 857 1912 891
rect 1946 857 1955 891
rect 1903 819 1955 857
rect 1903 785 1912 819
rect 1946 785 1955 819
rect 1903 747 1955 785
rect 1903 713 1912 747
rect 1946 713 1955 747
rect 1903 675 1955 713
rect 1903 641 1912 675
rect 1946 641 1955 675
rect 1903 639 1955 641
rect 1903 575 1912 587
rect 1946 575 1955 587
rect 1903 511 1912 523
rect 1946 511 1955 523
rect 1903 447 1912 459
rect 1946 447 1955 459
rect 1903 387 1955 395
rect 1903 383 1912 387
rect 1946 383 1955 387
rect 1903 319 1955 331
rect 1903 255 1955 267
rect 1903 197 1955 203
rect 2198 1179 2257 1191
rect 2198 1145 2204 1179
rect 2238 1145 2257 1179
rect 2198 1107 2257 1145
rect 2198 1073 2204 1107
rect 2238 1073 2257 1107
rect 2198 1035 2257 1073
rect 2198 1001 2204 1035
rect 2238 1001 2257 1035
rect 2198 963 2257 1001
rect 2198 929 2204 963
rect 2238 929 2257 963
rect 2198 891 2257 929
rect 2198 857 2204 891
rect 2238 857 2257 891
rect 2198 819 2257 857
rect 2198 785 2204 819
rect 2238 785 2257 819
rect 2198 747 2257 785
rect 2198 713 2204 747
rect 2238 713 2257 747
rect 2198 675 2257 713
rect 2198 641 2204 675
rect 2238 641 2257 675
rect 2198 603 2257 641
rect 2198 569 2204 603
rect 2238 569 2257 603
rect 2198 531 2257 569
rect 2198 497 2204 531
rect 2238 497 2257 531
rect 2198 459 2257 497
rect 2198 425 2204 459
rect 2238 425 2257 459
rect 2198 387 2257 425
rect 2198 353 2204 387
rect 2238 353 2257 387
rect 2198 315 2257 353
rect 2198 281 2204 315
rect 2238 281 2257 315
rect 2198 243 2257 281
rect 2198 209 2204 243
rect 2238 209 2257 243
rect 2198 197 2257 209
rect 381 125 1917 137
rect 381 19 412 125
rect 1886 19 1917 125
rect 381 0 1917 19
<< via1 >>
rect 343 603 395 639
rect 343 587 352 603
rect 352 587 386 603
rect 386 587 395 603
rect 343 569 352 575
rect 352 569 386 575
rect 386 569 395 575
rect 343 531 395 569
rect 343 523 352 531
rect 352 523 386 531
rect 386 523 395 531
rect 343 497 352 511
rect 352 497 386 511
rect 386 497 395 511
rect 343 459 395 497
rect 343 425 352 447
rect 352 425 386 447
rect 386 425 395 447
rect 343 395 395 425
rect 343 353 352 383
rect 352 353 386 383
rect 386 353 395 383
rect 343 331 395 353
rect 343 315 395 319
rect 343 281 352 315
rect 352 281 386 315
rect 386 281 395 315
rect 343 267 395 281
rect 343 243 395 255
rect 343 209 352 243
rect 352 209 386 243
rect 386 209 395 243
rect 343 203 395 209
rect 499 1179 551 1185
rect 499 1145 508 1179
rect 508 1145 542 1179
rect 542 1145 551 1179
rect 499 1133 551 1145
rect 499 1107 551 1121
rect 499 1073 508 1107
rect 508 1073 542 1107
rect 542 1073 551 1107
rect 499 1069 551 1073
rect 499 1035 551 1057
rect 499 1005 508 1035
rect 508 1005 542 1035
rect 542 1005 551 1035
rect 499 963 551 993
rect 499 941 508 963
rect 508 941 542 963
rect 542 941 551 963
rect 499 891 551 929
rect 499 877 508 891
rect 508 877 542 891
rect 542 877 551 891
rect 499 857 508 865
rect 508 857 542 865
rect 542 857 551 865
rect 499 819 551 857
rect 499 813 508 819
rect 508 813 542 819
rect 542 813 551 819
rect 499 785 508 801
rect 508 785 542 801
rect 542 785 551 801
rect 499 749 551 785
rect 655 603 707 639
rect 655 587 664 603
rect 664 587 698 603
rect 698 587 707 603
rect 655 569 664 575
rect 664 569 698 575
rect 698 569 707 575
rect 655 531 707 569
rect 655 523 664 531
rect 664 523 698 531
rect 698 523 707 531
rect 655 497 664 511
rect 664 497 698 511
rect 698 497 707 511
rect 655 459 707 497
rect 655 425 664 447
rect 664 425 698 447
rect 698 425 707 447
rect 655 395 707 425
rect 655 353 664 383
rect 664 353 698 383
rect 698 353 707 383
rect 655 331 707 353
rect 655 315 707 319
rect 655 281 664 315
rect 664 281 698 315
rect 698 281 707 315
rect 655 267 707 281
rect 655 243 707 255
rect 655 209 664 243
rect 664 209 698 243
rect 698 209 707 243
rect 655 203 707 209
rect 811 1179 863 1185
rect 811 1145 820 1179
rect 820 1145 854 1179
rect 854 1145 863 1179
rect 811 1133 863 1145
rect 811 1107 863 1121
rect 811 1073 820 1107
rect 820 1073 854 1107
rect 854 1073 863 1107
rect 811 1069 863 1073
rect 811 1035 863 1057
rect 811 1005 820 1035
rect 820 1005 854 1035
rect 854 1005 863 1035
rect 811 963 863 993
rect 811 941 820 963
rect 820 941 854 963
rect 854 941 863 963
rect 811 891 863 929
rect 811 877 820 891
rect 820 877 854 891
rect 854 877 863 891
rect 811 857 820 865
rect 820 857 854 865
rect 854 857 863 865
rect 811 819 863 857
rect 811 813 820 819
rect 820 813 854 819
rect 854 813 863 819
rect 811 785 820 801
rect 820 785 854 801
rect 854 785 863 801
rect 811 749 863 785
rect 967 603 1019 639
rect 967 587 976 603
rect 976 587 1010 603
rect 1010 587 1019 603
rect 967 569 976 575
rect 976 569 1010 575
rect 1010 569 1019 575
rect 967 531 1019 569
rect 967 523 976 531
rect 976 523 1010 531
rect 1010 523 1019 531
rect 967 497 976 511
rect 976 497 1010 511
rect 1010 497 1019 511
rect 967 459 1019 497
rect 967 425 976 447
rect 976 425 1010 447
rect 1010 425 1019 447
rect 967 395 1019 425
rect 967 353 976 383
rect 976 353 1010 383
rect 1010 353 1019 383
rect 967 331 1019 353
rect 967 315 1019 319
rect 967 281 976 315
rect 976 281 1010 315
rect 1010 281 1019 315
rect 967 267 1019 281
rect 967 243 1019 255
rect 967 209 976 243
rect 976 209 1010 243
rect 1010 209 1019 243
rect 967 203 1019 209
rect 1123 1179 1175 1185
rect 1123 1145 1132 1179
rect 1132 1145 1166 1179
rect 1166 1145 1175 1179
rect 1123 1133 1175 1145
rect 1123 1107 1175 1121
rect 1123 1073 1132 1107
rect 1132 1073 1166 1107
rect 1166 1073 1175 1107
rect 1123 1069 1175 1073
rect 1123 1035 1175 1057
rect 1123 1005 1132 1035
rect 1132 1005 1166 1035
rect 1166 1005 1175 1035
rect 1123 963 1175 993
rect 1123 941 1132 963
rect 1132 941 1166 963
rect 1166 941 1175 963
rect 1123 891 1175 929
rect 1123 877 1132 891
rect 1132 877 1166 891
rect 1166 877 1175 891
rect 1123 857 1132 865
rect 1132 857 1166 865
rect 1166 857 1175 865
rect 1123 819 1175 857
rect 1123 813 1132 819
rect 1132 813 1166 819
rect 1166 813 1175 819
rect 1123 785 1132 801
rect 1132 785 1166 801
rect 1166 785 1175 801
rect 1123 749 1175 785
rect 1279 603 1331 639
rect 1279 587 1288 603
rect 1288 587 1322 603
rect 1322 587 1331 603
rect 1279 569 1288 575
rect 1288 569 1322 575
rect 1322 569 1331 575
rect 1279 531 1331 569
rect 1279 523 1288 531
rect 1288 523 1322 531
rect 1322 523 1331 531
rect 1279 497 1288 511
rect 1288 497 1322 511
rect 1322 497 1331 511
rect 1279 459 1331 497
rect 1279 425 1288 447
rect 1288 425 1322 447
rect 1322 425 1331 447
rect 1279 395 1331 425
rect 1279 353 1288 383
rect 1288 353 1322 383
rect 1322 353 1331 383
rect 1279 331 1331 353
rect 1279 315 1331 319
rect 1279 281 1288 315
rect 1288 281 1322 315
rect 1322 281 1331 315
rect 1279 267 1331 281
rect 1279 243 1331 255
rect 1279 209 1288 243
rect 1288 209 1322 243
rect 1322 209 1331 243
rect 1279 203 1331 209
rect 1435 1179 1487 1185
rect 1435 1145 1444 1179
rect 1444 1145 1478 1179
rect 1478 1145 1487 1179
rect 1435 1133 1487 1145
rect 1435 1107 1487 1121
rect 1435 1073 1444 1107
rect 1444 1073 1478 1107
rect 1478 1073 1487 1107
rect 1435 1069 1487 1073
rect 1435 1035 1487 1057
rect 1435 1005 1444 1035
rect 1444 1005 1478 1035
rect 1478 1005 1487 1035
rect 1435 963 1487 993
rect 1435 941 1444 963
rect 1444 941 1478 963
rect 1478 941 1487 963
rect 1435 891 1487 929
rect 1435 877 1444 891
rect 1444 877 1478 891
rect 1478 877 1487 891
rect 1435 857 1444 865
rect 1444 857 1478 865
rect 1478 857 1487 865
rect 1435 819 1487 857
rect 1435 813 1444 819
rect 1444 813 1478 819
rect 1478 813 1487 819
rect 1435 785 1444 801
rect 1444 785 1478 801
rect 1478 785 1487 801
rect 1435 749 1487 785
rect 1591 603 1643 639
rect 1591 587 1600 603
rect 1600 587 1634 603
rect 1634 587 1643 603
rect 1591 569 1600 575
rect 1600 569 1634 575
rect 1634 569 1643 575
rect 1591 531 1643 569
rect 1591 523 1600 531
rect 1600 523 1634 531
rect 1634 523 1643 531
rect 1591 497 1600 511
rect 1600 497 1634 511
rect 1634 497 1643 511
rect 1591 459 1643 497
rect 1591 425 1600 447
rect 1600 425 1634 447
rect 1634 425 1643 447
rect 1591 395 1643 425
rect 1591 353 1600 383
rect 1600 353 1634 383
rect 1634 353 1643 383
rect 1591 331 1643 353
rect 1591 315 1643 319
rect 1591 281 1600 315
rect 1600 281 1634 315
rect 1634 281 1643 315
rect 1591 267 1643 281
rect 1591 243 1643 255
rect 1591 209 1600 243
rect 1600 209 1634 243
rect 1634 209 1643 243
rect 1591 203 1643 209
rect 1747 1179 1799 1185
rect 1747 1145 1756 1179
rect 1756 1145 1790 1179
rect 1790 1145 1799 1179
rect 1747 1133 1799 1145
rect 1747 1107 1799 1121
rect 1747 1073 1756 1107
rect 1756 1073 1790 1107
rect 1790 1073 1799 1107
rect 1747 1069 1799 1073
rect 1747 1035 1799 1057
rect 1747 1005 1756 1035
rect 1756 1005 1790 1035
rect 1790 1005 1799 1035
rect 1747 963 1799 993
rect 1747 941 1756 963
rect 1756 941 1790 963
rect 1790 941 1799 963
rect 1747 891 1799 929
rect 1747 877 1756 891
rect 1756 877 1790 891
rect 1790 877 1799 891
rect 1747 857 1756 865
rect 1756 857 1790 865
rect 1790 857 1799 865
rect 1747 819 1799 857
rect 1747 813 1756 819
rect 1756 813 1790 819
rect 1790 813 1799 819
rect 1747 785 1756 801
rect 1756 785 1790 801
rect 1790 785 1799 801
rect 1747 749 1799 785
rect 1903 603 1955 639
rect 1903 587 1912 603
rect 1912 587 1946 603
rect 1946 587 1955 603
rect 1903 569 1912 575
rect 1912 569 1946 575
rect 1946 569 1955 575
rect 1903 531 1955 569
rect 1903 523 1912 531
rect 1912 523 1946 531
rect 1946 523 1955 531
rect 1903 497 1912 511
rect 1912 497 1946 511
rect 1946 497 1955 511
rect 1903 459 1955 497
rect 1903 425 1912 447
rect 1912 425 1946 447
rect 1946 425 1955 447
rect 1903 395 1955 425
rect 1903 353 1912 383
rect 1912 353 1946 383
rect 1946 353 1955 383
rect 1903 331 1955 353
rect 1903 315 1955 319
rect 1903 281 1912 315
rect 1912 281 1946 315
rect 1946 281 1955 315
rect 1903 267 1955 281
rect 1903 243 1955 255
rect 1903 209 1912 243
rect 1912 209 1946 243
rect 1946 209 1955 243
rect 1903 203 1955 209
<< metal2 >>
rect 14 1185 2284 1191
rect 14 1133 499 1185
rect 551 1133 811 1185
rect 863 1133 1123 1185
rect 1175 1133 1435 1185
rect 1487 1133 1747 1185
rect 1799 1133 2284 1185
rect 14 1121 2284 1133
rect 14 1069 499 1121
rect 551 1069 811 1121
rect 863 1069 1123 1121
rect 1175 1069 1435 1121
rect 1487 1069 1747 1121
rect 1799 1069 2284 1121
rect 14 1057 2284 1069
rect 14 1005 499 1057
rect 551 1005 811 1057
rect 863 1005 1123 1057
rect 1175 1005 1435 1057
rect 1487 1005 1747 1057
rect 1799 1005 2284 1057
rect 14 993 2284 1005
rect 14 941 499 993
rect 551 941 811 993
rect 863 941 1123 993
rect 1175 941 1435 993
rect 1487 941 1747 993
rect 1799 941 2284 993
rect 14 929 2284 941
rect 14 877 499 929
rect 551 877 811 929
rect 863 877 1123 929
rect 1175 877 1435 929
rect 1487 877 1747 929
rect 1799 877 2284 929
rect 14 865 2284 877
rect 14 813 499 865
rect 551 813 811 865
rect 863 813 1123 865
rect 1175 813 1435 865
rect 1487 813 1747 865
rect 1799 813 2284 865
rect 14 801 2284 813
rect 14 749 499 801
rect 551 749 811 801
rect 863 749 1123 801
rect 1175 749 1435 801
rect 1487 749 1747 801
rect 1799 749 2284 801
rect 14 719 2284 749
rect 14 639 2284 669
rect 14 587 343 639
rect 395 587 655 639
rect 707 587 967 639
rect 1019 587 1279 639
rect 1331 587 1591 639
rect 1643 587 1903 639
rect 1955 587 2284 639
rect 14 575 2284 587
rect 14 523 343 575
rect 395 523 655 575
rect 707 523 967 575
rect 1019 523 1279 575
rect 1331 523 1591 575
rect 1643 523 1903 575
rect 1955 523 2284 575
rect 14 511 2284 523
rect 14 459 343 511
rect 395 459 655 511
rect 707 459 967 511
rect 1019 459 1279 511
rect 1331 459 1591 511
rect 1643 459 1903 511
rect 1955 459 2284 511
rect 14 447 2284 459
rect 14 395 343 447
rect 395 395 655 447
rect 707 395 967 447
rect 1019 395 1279 447
rect 1331 395 1591 447
rect 1643 395 1903 447
rect 1955 395 2284 447
rect 14 383 2284 395
rect 14 331 343 383
rect 395 331 655 383
rect 707 331 967 383
rect 1019 331 1279 383
rect 1331 331 1591 383
rect 1643 331 1903 383
rect 1955 331 2284 383
rect 14 319 2284 331
rect 14 267 343 319
rect 395 267 655 319
rect 707 267 967 319
rect 1019 267 1279 319
rect 1331 267 1591 319
rect 1643 267 1903 319
rect 1955 267 2284 319
rect 14 255 2284 267
rect 14 203 343 255
rect 395 203 655 255
rect 707 203 967 255
rect 1019 203 1279 255
rect 1331 203 1591 255
rect 1643 203 1903 255
rect 1955 203 2284 255
rect 14 197 2284 203
<< labels >>
flabel comment s 2005 687 2005 687 0 FreeSans 400 90 0 0 dummy_poly
flabel comment s 283 660 283 660 0 FreeSans 400 90 0 0 dummy_poly
flabel metal1 s 1098 85 1195 120 0 FreeSans 200 0 0 0 GATE
port 3 nsew
flabel metal1 s 2198 679 2257 709 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal1 s 41 675 100 705 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal2 s 25 442 128 488 0 FreeSans 200 0 0 0 SOURCE
port 4 nsew
flabel metal2 s 25 991 137 1048 0 FreeSans 200 0 0 0 DRAIN
port 5 nsew
<< properties >>
string GDS_END 8608414
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8555078
<< end >>
