magic
tech sky130B
magscale 1 2
timestamp 1688980957
use sky130_fd_pr__nfet_01v8__example_55959141808571  sky130_fd_pr__nfet_01v8__example_55959141808571_0
timestamp 1688980957
transform 1 0 119 0 1 36
box -1 0 297 1
use sky130_fd_pr__pfet_01v8__example_55959141808441  sky130_fd_pr__pfet_01v8__example_55959141808441_0
timestamp 1688980957
transform 1 0 119 0 1 350
box -1 0 297 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1688980957
transform -1 0 205 0 -1 302
box 0 0 1 1
<< properties >>
string GDS_END 8157834
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8155234
<< end >>
