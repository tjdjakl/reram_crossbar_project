magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 157 439 203
rect 1538 157 2006 203
rect 1 21 2006 157
rect 30 -17 64 21
<< locali >>
rect 103 317 169 489
rect 287 390 329 493
rect 280 356 329 390
rect 280 317 314 356
rect 17 283 314 317
rect 650 314 868 348
rect 17 181 87 283
rect 17 147 305 181
rect 103 51 169 147
rect 271 97 305 147
rect 650 255 684 314
rect 610 221 684 255
rect 834 250 868 314
rect 1319 337 1369 391
rect 1044 303 1369 337
rect 1044 287 1116 303
rect 1044 250 1078 287
rect 1319 271 1369 303
rect 1664 393 1698 493
rect 1664 359 1714 393
rect 834 193 1078 250
rect 1680 317 1714 359
rect 1832 317 1898 485
rect 1680 283 2007 317
rect 271 63 337 97
rect 1940 181 2007 283
rect 1680 147 2007 181
rect 1680 97 1730 147
rect 1664 51 1730 97
rect 1832 54 1898 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 35 359 69 527
rect 203 359 237 527
rect 363 455 429 527
rect 547 416 634 493
rect 428 382 634 416
rect 668 421 702 493
rect 736 455 802 527
rect 836 421 883 493
rect 668 387 883 421
rect 924 383 990 527
rect 1024 421 1058 493
rect 1092 455 1158 527
rect 1192 421 1226 493
rect 1282 425 1522 493
rect 1563 455 1629 527
rect 1024 387 1226 421
rect 1488 421 1522 425
rect 428 333 462 382
rect 355 320 462 333
rect 348 299 462 320
rect 496 323 616 338
rect 348 286 389 299
rect 496 289 582 323
rect 348 249 382 286
rect 121 215 382 249
rect 35 17 69 113
rect 203 17 237 113
rect 348 165 382 215
rect 416 255 468 265
rect 416 221 490 255
rect 524 221 536 255
rect 722 255 800 272
rect 722 221 766 255
rect 416 199 536 221
rect 722 206 800 221
rect 916 323 999 349
rect 1488 387 1621 421
rect 916 289 954 323
rect 988 289 999 323
rect 916 287 999 289
rect 1415 323 1552 347
rect 1415 289 1506 323
rect 1540 289 1552 323
rect 1587 328 1621 387
rect 1748 359 1782 527
rect 1587 294 1645 328
rect 1129 221 1138 255
rect 1172 221 1201 255
rect 1129 191 1201 221
rect 1235 191 1372 225
rect 1406 221 1414 255
rect 1448 221 1577 255
rect 1406 199 1577 221
rect 1611 249 1645 294
rect 1932 359 1966 527
rect 1611 215 1889 249
rect 570 165 618 187
rect 348 131 618 165
rect 371 17 437 93
rect 474 51 618 131
rect 668 123 870 157
rect 668 51 702 123
rect 736 17 802 89
rect 836 51 870 123
rect 1024 123 1226 157
rect 1269 153 1372 191
rect 1611 165 1645 215
rect 924 17 990 98
rect 1024 51 1058 123
rect 1092 17 1158 89
rect 1192 51 1226 123
rect 1461 131 1645 165
rect 1293 101 1327 119
rect 1461 101 1495 131
rect 1293 51 1495 101
rect 1541 17 1607 89
rect 1764 17 1798 113
rect 1932 17 1966 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 582 289 616 323
rect 490 221 524 255
rect 766 221 800 255
rect 954 289 988 323
rect 1506 289 1540 323
rect 1138 221 1172 255
rect 1414 221 1448 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 570 323 628 329
rect 570 289 582 323
rect 616 320 628 323
rect 942 323 1000 329
rect 942 320 954 323
rect 616 292 954 320
rect 616 289 628 292
rect 570 283 628 289
rect 942 289 954 292
rect 988 320 1000 323
rect 1494 323 1552 329
rect 1494 320 1506 323
rect 988 292 1506 320
rect 988 289 1000 292
rect 942 283 1000 289
rect 1494 289 1506 292
rect 1540 289 1552 323
rect 1494 283 1552 289
rect 478 255 536 261
rect 478 221 490 255
rect 524 252 536 255
rect 754 255 812 261
rect 754 252 766 255
rect 524 224 766 252
rect 524 221 536 224
rect 478 215 536 221
rect 754 221 766 224
rect 800 252 812 255
rect 1126 255 1184 261
rect 1126 252 1138 255
rect 800 224 1138 252
rect 800 221 812 224
rect 754 215 812 221
rect 1126 221 1138 224
rect 1172 252 1184 255
rect 1402 255 1460 261
rect 1402 252 1414 255
rect 1172 224 1414 252
rect 1172 221 1184 224
rect 1126 215 1184 221
rect 1402 221 1414 224
rect 1448 221 1460 255
rect 1402 215 1460 221
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< obsm1 >>
rect 570 184 628 193
rect 1310 184 1368 193
rect 570 156 1368 184
rect 570 147 628 156
rect 1310 147 1368 156
<< labels >>
rlabel metal1 s 1402 215 1460 224 6 A
port 1 nsew signal input
rlabel metal1 s 1126 215 1184 224 6 A
port 1 nsew signal input
rlabel metal1 s 754 215 812 224 6 A
port 1 nsew signal input
rlabel metal1 s 478 215 536 224 6 A
port 1 nsew signal input
rlabel metal1 s 478 224 1460 252 6 A
port 1 nsew signal input
rlabel metal1 s 1402 252 1460 261 6 A
port 1 nsew signal input
rlabel metal1 s 1126 252 1184 261 6 A
port 1 nsew signal input
rlabel metal1 s 754 252 812 261 6 A
port 1 nsew signal input
rlabel metal1 s 478 252 536 261 6 A
port 1 nsew signal input
rlabel metal1 s 1494 283 1552 292 6 B
port 2 nsew signal input
rlabel metal1 s 942 283 1000 292 6 B
port 2 nsew signal input
rlabel metal1 s 570 283 628 292 6 B
port 2 nsew signal input
rlabel metal1 s 570 292 1552 320 6 B
port 2 nsew signal input
rlabel metal1 s 1494 320 1552 329 6 B
port 2 nsew signal input
rlabel metal1 s 942 320 1000 329 6 B
port 2 nsew signal input
rlabel metal1 s 570 320 628 329 6 B
port 2 nsew signal input
rlabel locali s 834 193 1078 250 6 CIN
port 3 nsew signal input
rlabel locali s 1319 271 1369 303 6 CIN
port 3 nsew signal input
rlabel locali s 1044 250 1078 287 6 CIN
port 3 nsew signal input
rlabel locali s 1044 287 1116 303 6 CIN
port 3 nsew signal input
rlabel locali s 1044 303 1369 337 6 CIN
port 3 nsew signal input
rlabel locali s 834 250 868 314 6 CIN
port 3 nsew signal input
rlabel locali s 610 221 684 255 6 CIN
port 3 nsew signal input
rlabel locali s 650 255 684 314 6 CIN
port 3 nsew signal input
rlabel locali s 1319 337 1369 391 6 CIN
port 3 nsew signal input
rlabel locali s 650 314 868 348 6 CIN
port 3 nsew signal input
rlabel metal1 s 0 -48 2024 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 2006 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1538 157 2006 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 157 439 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 271 63 337 97 6 COUT
port 8 nsew signal output
rlabel locali s 271 97 305 147 6 COUT
port 8 nsew signal output
rlabel locali s 103 51 169 147 6 COUT
port 8 nsew signal output
rlabel locali s 17 147 305 181 6 COUT
port 8 nsew signal output
rlabel locali s 17 181 87 283 6 COUT
port 8 nsew signal output
rlabel locali s 17 283 314 317 6 COUT
port 8 nsew signal output
rlabel locali s 280 317 314 356 6 COUT
port 8 nsew signal output
rlabel locali s 280 356 329 390 6 COUT
port 8 nsew signal output
rlabel locali s 287 390 329 493 6 COUT
port 8 nsew signal output
rlabel locali s 103 317 169 489 6 COUT
port 8 nsew signal output
rlabel locali s 1832 54 1898 147 6 SUM
port 9 nsew signal output
rlabel locali s 1664 51 1730 97 6 SUM
port 9 nsew signal output
rlabel locali s 1680 97 1730 147 6 SUM
port 9 nsew signal output
rlabel locali s 1680 147 2007 181 6 SUM
port 9 nsew signal output
rlabel locali s 1940 181 2007 283 6 SUM
port 9 nsew signal output
rlabel locali s 1680 283 2007 317 6 SUM
port 9 nsew signal output
rlabel locali s 1832 317 1898 485 6 SUM
port 9 nsew signal output
rlabel locali s 1680 317 1714 359 6 SUM
port 9 nsew signal output
rlabel locali s 1664 359 1714 393 6 SUM
port 9 nsew signal output
rlabel locali s 1664 393 1698 493 6 SUM
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2024 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2093974
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2078288
<< end >>
