magic
tech sky130B
magscale 1 2
timestamp 1700624956
<< locali >>
rect 214 2496 930 2536
rect 214 2364 446 2496
rect 904 2364 930 2496
rect 214 2212 930 2364
rect 214 2156 342 2212
rect 214 2034 356 2156
rect 214 1504 342 2034
rect 802 1504 930 2212
rect 214 702 342 1252
rect 758 702 932 1252
rect 214 600 932 702
rect 214 468 448 600
rect 906 468 932 600
rect 214 420 932 468
<< viali >>
rect 446 2364 904 2496
rect 448 468 906 600
<< metal1 >>
rect 214 2496 930 2536
rect 214 2364 446 2496
rect 904 2364 930 2496
rect 214 2226 930 2364
rect 128 2110 328 2162
rect 128 2064 602 2110
rect 128 1962 328 2064
rect 128 1402 328 1466
rect 454 1402 496 1944
rect 550 1640 594 2064
rect 128 1334 496 1402
rect 128 1266 328 1334
rect 454 958 496 1334
rect 648 1402 690 1948
rect 816 1402 1016 1466
rect 648 1334 1016 1402
rect 126 860 326 954
rect 550 860 592 1112
rect 648 962 690 1334
rect 816 1266 1016 1334
rect 126 814 544 860
rect 126 754 326 814
rect 214 600 932 640
rect 214 468 448 600
rect 906 468 932 600
rect 214 420 932 468
use sky130_fd_pr__nfet_g5v0d10v5_6XHARQ  XM1
timestamp 1700618825
transform 1 0 572 0 1 967
box -278 -333 278 333
use sky130_fd_pr__pfet_g5v0d10v5_7EBZY6  XM2
timestamp 1700618825
transform 1 0 572 0 1 1873
box -308 -447 308 447
<< labels >>
flabel metal1 228 2328 428 2528 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 230 432 430 632 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 128 1266 328 1466 0 FreeSans 256 0 0 0 In
port 1 nsew
flabel metal1 816 1266 1016 1466 0 FreeSans 256 0 0 0 Out
port 0 nsew
flabel metal1 128 1962 328 2162 0 FreeSans 256 0 0 0 SP
port 2 nsew
flabel metal1 126 754 326 954 0 FreeSans 256 0 0 0 SN
port 5 nsew
<< end >>
