magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< pwell >>
rect -13 -26 73 1246
rect 257 572 278 621
rect 467 -26 553 1246
<< locali >>
rect 13 0 47 1220
rect 493 0 527 1220
<< metal1 >>
rect 14 1213 526 1220
rect 14 1161 44 1213
rect 96 1161 284 1213
rect 336 1161 364 1213
rect 416 1161 444 1213
rect 496 1161 526 1213
rect 14 1154 526 1161
rect 14 126 46 1154
rect 74 66 106 1094
rect 134 126 166 1154
rect 194 66 226 1094
rect 254 126 286 1154
rect 314 66 346 1094
rect 374 126 406 1154
rect 434 66 466 1094
rect 494 126 526 1154
rect 60 59 480 66
rect 60 7 84 59
rect 136 7 164 59
rect 216 7 244 59
rect 296 7 324 59
rect 376 7 404 59
rect 456 7 480 59
rect 60 0 480 7
<< via1 >>
rect 44 1161 96 1213
rect 284 1161 336 1213
rect 364 1161 416 1213
rect 444 1161 496 1213
rect 84 7 136 59
rect 164 7 216 59
rect 244 7 296 59
rect 324 7 376 59
rect 404 7 456 59
<< metal2 >>
rect 14 1215 166 1220
rect 14 1159 42 1215
rect 98 1159 166 1215
rect 14 1154 166 1159
rect 14 126 46 1154
rect 74 66 106 1094
rect 134 126 166 1154
rect 194 66 226 1220
rect 254 1215 526 1220
rect 254 1159 282 1215
rect 338 1159 362 1215
rect 418 1159 442 1215
rect 498 1159 526 1215
rect 254 1154 526 1159
rect 254 126 286 1154
rect 314 66 346 1094
rect 374 126 406 1154
rect 434 66 466 1094
rect 494 126 526 1154
rect 60 61 480 66
rect 60 5 82 61
rect 138 5 162 61
rect 218 5 242 61
rect 298 5 322 61
rect 378 5 402 61
rect 458 5 480 61
rect 60 0 480 5
<< via2 >>
rect 42 1213 98 1215
rect 42 1161 44 1213
rect 44 1161 96 1213
rect 96 1161 98 1213
rect 42 1159 98 1161
rect 282 1213 338 1215
rect 282 1161 284 1213
rect 284 1161 336 1213
rect 336 1161 338 1213
rect 282 1159 338 1161
rect 362 1213 418 1215
rect 362 1161 364 1213
rect 364 1161 416 1213
rect 416 1161 418 1213
rect 362 1159 418 1161
rect 442 1213 498 1215
rect 442 1161 444 1213
rect 444 1161 496 1213
rect 496 1161 498 1213
rect 442 1159 498 1161
rect 82 59 138 61
rect 82 7 84 59
rect 84 7 136 59
rect 136 7 138 59
rect 82 5 138 7
rect 162 59 218 61
rect 162 7 164 59
rect 164 7 216 59
rect 216 7 218 59
rect 162 5 218 7
rect 242 59 298 61
rect 242 7 244 59
rect 244 7 296 59
rect 296 7 298 59
rect 242 5 298 7
rect 322 59 378 61
rect 322 7 324 59
rect 324 7 376 59
rect 376 7 378 59
rect 322 5 378 7
rect 402 59 458 61
rect 402 7 404 59
rect 404 7 456 59
rect 456 7 458 59
rect 402 5 458 7
<< metal3 >>
rect 0 1219 540 1220
rect 0 1155 38 1219
rect 102 1155 118 1219
rect 182 1155 198 1219
rect 262 1155 278 1219
rect 342 1155 358 1219
rect 422 1155 438 1219
rect 502 1155 540 1219
rect 0 1154 540 1155
rect 0 126 60 1154
rect 120 66 180 1094
rect 240 126 300 1154
rect 360 66 420 1094
rect 480 126 540 1154
rect 60 65 480 66
rect 60 1 78 65
rect 142 1 158 65
rect 222 1 238 65
rect 302 1 318 65
rect 382 1 398 65
rect 462 1 480 65
rect 60 0 480 1
<< via3 >>
rect 38 1215 102 1219
rect 38 1159 42 1215
rect 42 1159 98 1215
rect 98 1159 102 1215
rect 38 1155 102 1159
rect 118 1155 182 1219
rect 198 1155 262 1219
rect 278 1215 342 1219
rect 278 1159 282 1215
rect 282 1159 338 1215
rect 338 1159 342 1215
rect 278 1155 342 1159
rect 358 1215 422 1219
rect 358 1159 362 1215
rect 362 1159 418 1215
rect 418 1159 422 1215
rect 358 1155 422 1159
rect 438 1215 502 1219
rect 438 1159 442 1215
rect 442 1159 498 1215
rect 498 1159 502 1215
rect 438 1155 502 1159
rect 78 61 142 65
rect 78 5 82 61
rect 82 5 138 61
rect 138 5 142 61
rect 78 1 142 5
rect 158 61 222 65
rect 158 5 162 61
rect 162 5 218 61
rect 218 5 222 61
rect 158 1 222 5
rect 238 61 302 65
rect 238 5 242 61
rect 242 5 298 61
rect 298 5 302 61
rect 238 1 302 5
rect 318 61 382 65
rect 318 5 322 61
rect 322 5 378 61
rect 378 5 382 61
rect 318 1 382 5
rect 398 61 462 65
rect 398 5 402 61
rect 402 5 458 61
rect 458 5 462 61
rect 398 1 462 5
<< metal4 >>
rect 0 1219 540 1220
rect 0 1155 38 1219
rect 102 1155 118 1219
rect 182 1155 198 1219
rect 262 1155 278 1219
rect 342 1155 358 1219
rect 422 1155 438 1219
rect 502 1155 540 1219
rect 0 1154 540 1155
rect 0 126 60 1154
rect 120 66 180 1094
rect 240 126 300 1154
rect 360 66 420 1094
rect 480 126 540 1154
rect 60 65 480 66
rect 60 1 78 65
rect 142 1 158 65
rect 222 1 238 65
rect 302 1 318 65
rect 382 1 398 65
rect 462 1 480 65
rect 60 0 480 1
<< labels >>
flabel metal2 s 140 270 159 290 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 287 21 323 57 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 257 572 278 621 0 FreeSans 400 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 10464
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 4272
string path 1.500 0.825 12.000 0.825 
<< end >>
