magic
tech sky130B
magscale 1 2
timestamp 1688980957
use sky130_fd_pr__hvdfl1sd2__example_55959141808316  sky130_fd_pr__hvdfl1sd2__example_55959141808316_0
timestamp 1688980957
transform 1 0 800 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808137  sky130_fd_pr__hvdfl1sd__example_55959141808137_0
timestamp 1688980957
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808137  sky130_fd_pr__hvdfl1sd__example_55959141808137_1
timestamp 1688980957
transform 1 0 1656 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 37016432
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37014860
<< end >>
