magic
tech sky130B
magscale 1 2
timestamp 1688980957
use sky130_fd_io__nfet_con_diff_wo_abt_270v2  sky130_fd_io__nfet_con_diff_wo_abt_270v2_0
timestamp 1688980957
transform -1 0 15088 0 -1 8404
box 0 423 15173 5493
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_0
timestamp 1688980957
transform 0 -1 12892 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_1
timestamp 1688980957
transform 0 -1 11458 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_2
timestamp 1688980957
transform 0 -1 10115 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_3
timestamp 1688980957
transform 0 -1 8635 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_4
timestamp 1688980957
transform 0 -1 6933 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_5
timestamp 1688980957
transform 0 -1 13322 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_6
timestamp 1688980957
transform 0 -1 10975 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_7
timestamp 1688980957
transform 0 -1 9495 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_8
timestamp 1688980957
transform 0 -1 12318 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_9
timestamp 1688980957
transform 0 -1 7793 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_10
timestamp 1688980957
transform 0 -1 1977 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_11
timestamp 1688980957
transform 0 -1 1694 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_12
timestamp 1688980957
transform 0 1 413 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_13
timestamp 1688980957
transform 0 1 896 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_0
timestamp 1688980957
transform 0 -1 11888 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_1
timestamp 1688980957
transform 0 -1 7363 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_2
timestamp 1688980957
transform 0 -1 10545 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_3
timestamp 1688980957
transform 0 -1 9065 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_4
timestamp 1688980957
transform 0 -1 13752 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_5
timestamp 1688980957
transform 0 -1 1390 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_6
timestamp 1688980957
transform 0 1 655 1 0 1584
box 0 0 1 1
use sky130_fd_pr__res_generic_po__example_5595914180838  sky130_fd_pr__res_generic_po__example_5595914180838_0
timestamp 1688980957
transform 1 0 336 0 1 9367
box 15 17 2025 18
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_0
timestamp 1688980957
transform -1 0 2461 0 -1 9417
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_1
timestamp 1688980957
transform 1 0 251 0 -1 9417
box 0 0 1 1
<< properties >>
string GDS_END 4473848
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 4438700
<< end >>
