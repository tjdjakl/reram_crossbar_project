magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< dnwell >>
rect -38 -38 1072 7440
<< nwell >>
rect -118 7319 168 7520
rect 782 7319 1119 7520
rect -118 7150 1119 7319
rect -118 168 168 7150
rect 782 168 1119 7150
rect -118 0 1119 168
rect 2 -76 948 0
<< pwell >>
rect 228 228 722 7090
<< mvnmos >>
rect 415 5956 535 6956
rect 415 4835 535 5835
rect 415 3714 535 4714
rect 415 2604 535 3604
rect 415 1483 535 2483
rect 415 362 535 1362
<< mvndiff >>
rect 362 6944 415 6956
rect 362 6910 370 6944
rect 404 6910 415 6944
rect 362 6876 415 6910
rect 362 6842 370 6876
rect 404 6842 415 6876
rect 362 6808 415 6842
rect 362 6774 370 6808
rect 404 6774 415 6808
rect 362 6740 415 6774
rect 362 6706 370 6740
rect 404 6706 415 6740
rect 362 6672 415 6706
rect 362 6638 370 6672
rect 404 6638 415 6672
rect 362 6604 415 6638
rect 362 6570 370 6604
rect 404 6570 415 6604
rect 362 6536 415 6570
rect 362 6502 370 6536
rect 404 6502 415 6536
rect 362 6468 415 6502
rect 362 6434 370 6468
rect 404 6434 415 6468
rect 362 6400 415 6434
rect 362 6366 370 6400
rect 404 6366 415 6400
rect 362 6332 415 6366
rect 362 6298 370 6332
rect 404 6298 415 6332
rect 362 6264 415 6298
rect 362 6230 370 6264
rect 404 6230 415 6264
rect 362 6196 415 6230
rect 362 6162 370 6196
rect 404 6162 415 6196
rect 362 6128 415 6162
rect 362 6094 370 6128
rect 404 6094 415 6128
rect 362 6060 415 6094
rect 362 6026 370 6060
rect 404 6026 415 6060
rect 362 5956 415 6026
rect 535 6944 588 6956
rect 535 6910 546 6944
rect 580 6910 588 6944
rect 535 6876 588 6910
rect 535 6842 546 6876
rect 580 6842 588 6876
rect 535 6808 588 6842
rect 535 6774 546 6808
rect 580 6774 588 6808
rect 535 6740 588 6774
rect 535 6706 546 6740
rect 580 6706 588 6740
rect 535 6672 588 6706
rect 535 6638 546 6672
rect 580 6638 588 6672
rect 535 6604 588 6638
rect 535 6570 546 6604
rect 580 6570 588 6604
rect 535 6536 588 6570
rect 535 6502 546 6536
rect 580 6502 588 6536
rect 535 6468 588 6502
rect 535 6434 546 6468
rect 580 6434 588 6468
rect 535 6400 588 6434
rect 535 6366 546 6400
rect 580 6366 588 6400
rect 535 6332 588 6366
rect 535 6298 546 6332
rect 580 6298 588 6332
rect 535 6264 588 6298
rect 535 6230 546 6264
rect 580 6230 588 6264
rect 535 6196 588 6230
rect 535 6162 546 6196
rect 580 6162 588 6196
rect 535 6128 588 6162
rect 535 6094 546 6128
rect 580 6094 588 6128
rect 535 6060 588 6094
rect 535 6026 546 6060
rect 580 6026 588 6060
rect 535 5956 588 6026
rect 362 5823 415 5835
rect 362 5789 370 5823
rect 404 5789 415 5823
rect 362 5755 415 5789
rect 362 5721 370 5755
rect 404 5721 415 5755
rect 362 5687 415 5721
rect 362 5653 370 5687
rect 404 5653 415 5687
rect 362 5619 415 5653
rect 362 5585 370 5619
rect 404 5585 415 5619
rect 362 5551 415 5585
rect 362 5517 370 5551
rect 404 5517 415 5551
rect 362 5483 415 5517
rect 362 5449 370 5483
rect 404 5449 415 5483
rect 362 5415 415 5449
rect 362 5381 370 5415
rect 404 5381 415 5415
rect 362 5347 415 5381
rect 362 5313 370 5347
rect 404 5313 415 5347
rect 362 5279 415 5313
rect 362 5245 370 5279
rect 404 5245 415 5279
rect 362 5211 415 5245
rect 362 5177 370 5211
rect 404 5177 415 5211
rect 362 5143 415 5177
rect 362 5109 370 5143
rect 404 5109 415 5143
rect 362 5075 415 5109
rect 362 5041 370 5075
rect 404 5041 415 5075
rect 362 5007 415 5041
rect 362 4973 370 5007
rect 404 4973 415 5007
rect 362 4939 415 4973
rect 362 4905 370 4939
rect 404 4905 415 4939
rect 362 4835 415 4905
rect 535 5823 588 5835
rect 535 5789 546 5823
rect 580 5789 588 5823
rect 535 5755 588 5789
rect 535 5721 546 5755
rect 580 5721 588 5755
rect 535 5687 588 5721
rect 535 5653 546 5687
rect 580 5653 588 5687
rect 535 5619 588 5653
rect 535 5585 546 5619
rect 580 5585 588 5619
rect 535 5551 588 5585
rect 535 5517 546 5551
rect 580 5517 588 5551
rect 535 5483 588 5517
rect 535 5449 546 5483
rect 580 5449 588 5483
rect 535 5415 588 5449
rect 535 5381 546 5415
rect 580 5381 588 5415
rect 535 5347 588 5381
rect 535 5313 546 5347
rect 580 5313 588 5347
rect 535 5279 588 5313
rect 535 5245 546 5279
rect 580 5245 588 5279
rect 535 5211 588 5245
rect 535 5177 546 5211
rect 580 5177 588 5211
rect 535 5143 588 5177
rect 535 5109 546 5143
rect 580 5109 588 5143
rect 535 5075 588 5109
rect 535 5041 546 5075
rect 580 5041 588 5075
rect 535 5007 588 5041
rect 535 4973 546 5007
rect 580 4973 588 5007
rect 535 4939 588 4973
rect 535 4905 546 4939
rect 580 4905 588 4939
rect 535 4835 588 4905
rect 362 4702 415 4714
rect 362 4668 370 4702
rect 404 4668 415 4702
rect 362 4634 415 4668
rect 362 4600 370 4634
rect 404 4600 415 4634
rect 362 4566 415 4600
rect 362 4532 370 4566
rect 404 4532 415 4566
rect 362 4498 415 4532
rect 362 4464 370 4498
rect 404 4464 415 4498
rect 362 4430 415 4464
rect 362 4396 370 4430
rect 404 4396 415 4430
rect 362 4362 415 4396
rect 362 4328 370 4362
rect 404 4328 415 4362
rect 362 4294 415 4328
rect 362 4260 370 4294
rect 404 4260 415 4294
rect 362 4226 415 4260
rect 362 4192 370 4226
rect 404 4192 415 4226
rect 362 4158 415 4192
rect 362 4124 370 4158
rect 404 4124 415 4158
rect 362 4090 415 4124
rect 362 4056 370 4090
rect 404 4056 415 4090
rect 362 4022 415 4056
rect 362 3988 370 4022
rect 404 3988 415 4022
rect 362 3954 415 3988
rect 362 3920 370 3954
rect 404 3920 415 3954
rect 362 3886 415 3920
rect 362 3852 370 3886
rect 404 3852 415 3886
rect 362 3818 415 3852
rect 362 3784 370 3818
rect 404 3784 415 3818
rect 362 3714 415 3784
rect 535 4702 588 4714
rect 535 4668 546 4702
rect 580 4668 588 4702
rect 535 4634 588 4668
rect 535 4600 546 4634
rect 580 4600 588 4634
rect 535 4566 588 4600
rect 535 4532 546 4566
rect 580 4532 588 4566
rect 535 4498 588 4532
rect 535 4464 546 4498
rect 580 4464 588 4498
rect 535 4430 588 4464
rect 535 4396 546 4430
rect 580 4396 588 4430
rect 535 4362 588 4396
rect 535 4328 546 4362
rect 580 4328 588 4362
rect 535 4294 588 4328
rect 535 4260 546 4294
rect 580 4260 588 4294
rect 535 4226 588 4260
rect 535 4192 546 4226
rect 580 4192 588 4226
rect 535 4158 588 4192
rect 535 4124 546 4158
rect 580 4124 588 4158
rect 535 4090 588 4124
rect 535 4056 546 4090
rect 580 4056 588 4090
rect 535 4022 588 4056
rect 535 3988 546 4022
rect 580 3988 588 4022
rect 535 3954 588 3988
rect 535 3920 546 3954
rect 580 3920 588 3954
rect 535 3886 588 3920
rect 535 3852 546 3886
rect 580 3852 588 3886
rect 535 3818 588 3852
rect 535 3784 546 3818
rect 580 3784 588 3818
rect 535 3714 588 3784
rect 362 3534 415 3604
rect 362 3500 370 3534
rect 404 3500 415 3534
rect 362 3466 415 3500
rect 362 3432 370 3466
rect 404 3432 415 3466
rect 362 3398 415 3432
rect 362 3364 370 3398
rect 404 3364 415 3398
rect 362 3330 415 3364
rect 362 3296 370 3330
rect 404 3296 415 3330
rect 362 3262 415 3296
rect 362 3228 370 3262
rect 404 3228 415 3262
rect 362 3194 415 3228
rect 362 3160 370 3194
rect 404 3160 415 3194
rect 362 3126 415 3160
rect 362 3092 370 3126
rect 404 3092 415 3126
rect 362 3058 415 3092
rect 362 3024 370 3058
rect 404 3024 415 3058
rect 362 2990 415 3024
rect 362 2956 370 2990
rect 404 2956 415 2990
rect 362 2922 415 2956
rect 362 2888 370 2922
rect 404 2888 415 2922
rect 362 2854 415 2888
rect 362 2820 370 2854
rect 404 2820 415 2854
rect 362 2786 415 2820
rect 362 2752 370 2786
rect 404 2752 415 2786
rect 362 2718 415 2752
rect 362 2684 370 2718
rect 404 2684 415 2718
rect 362 2650 415 2684
rect 362 2616 370 2650
rect 404 2616 415 2650
rect 362 2604 415 2616
rect 535 3534 588 3604
rect 535 3500 546 3534
rect 580 3500 588 3534
rect 535 3466 588 3500
rect 535 3432 546 3466
rect 580 3432 588 3466
rect 535 3398 588 3432
rect 535 3364 546 3398
rect 580 3364 588 3398
rect 535 3330 588 3364
rect 535 3296 546 3330
rect 580 3296 588 3330
rect 535 3262 588 3296
rect 535 3228 546 3262
rect 580 3228 588 3262
rect 535 3194 588 3228
rect 535 3160 546 3194
rect 580 3160 588 3194
rect 535 3126 588 3160
rect 535 3092 546 3126
rect 580 3092 588 3126
rect 535 3058 588 3092
rect 535 3024 546 3058
rect 580 3024 588 3058
rect 535 2990 588 3024
rect 535 2956 546 2990
rect 580 2956 588 2990
rect 535 2922 588 2956
rect 535 2888 546 2922
rect 580 2888 588 2922
rect 535 2854 588 2888
rect 535 2820 546 2854
rect 580 2820 588 2854
rect 535 2786 588 2820
rect 535 2752 546 2786
rect 580 2752 588 2786
rect 535 2718 588 2752
rect 535 2684 546 2718
rect 580 2684 588 2718
rect 535 2650 588 2684
rect 535 2616 546 2650
rect 580 2616 588 2650
rect 535 2604 588 2616
rect 362 2413 415 2483
rect 362 2379 370 2413
rect 404 2379 415 2413
rect 362 2345 415 2379
rect 362 2311 370 2345
rect 404 2311 415 2345
rect 362 2277 415 2311
rect 362 2243 370 2277
rect 404 2243 415 2277
rect 362 2209 415 2243
rect 362 2175 370 2209
rect 404 2175 415 2209
rect 362 2141 415 2175
rect 362 2107 370 2141
rect 404 2107 415 2141
rect 362 2073 415 2107
rect 362 2039 370 2073
rect 404 2039 415 2073
rect 362 2005 415 2039
rect 362 1971 370 2005
rect 404 1971 415 2005
rect 362 1937 415 1971
rect 362 1903 370 1937
rect 404 1903 415 1937
rect 362 1869 415 1903
rect 362 1835 370 1869
rect 404 1835 415 1869
rect 362 1801 415 1835
rect 362 1767 370 1801
rect 404 1767 415 1801
rect 362 1733 415 1767
rect 362 1699 370 1733
rect 404 1699 415 1733
rect 362 1665 415 1699
rect 362 1631 370 1665
rect 404 1631 415 1665
rect 362 1597 415 1631
rect 362 1563 370 1597
rect 404 1563 415 1597
rect 362 1529 415 1563
rect 362 1495 370 1529
rect 404 1495 415 1529
rect 362 1483 415 1495
rect 535 2413 588 2483
rect 535 2379 546 2413
rect 580 2379 588 2413
rect 535 2345 588 2379
rect 535 2311 546 2345
rect 580 2311 588 2345
rect 535 2277 588 2311
rect 535 2243 546 2277
rect 580 2243 588 2277
rect 535 2209 588 2243
rect 535 2175 546 2209
rect 580 2175 588 2209
rect 535 2141 588 2175
rect 535 2107 546 2141
rect 580 2107 588 2141
rect 535 2073 588 2107
rect 535 2039 546 2073
rect 580 2039 588 2073
rect 535 2005 588 2039
rect 535 1971 546 2005
rect 580 1971 588 2005
rect 535 1937 588 1971
rect 535 1903 546 1937
rect 580 1903 588 1937
rect 535 1869 588 1903
rect 535 1835 546 1869
rect 580 1835 588 1869
rect 535 1801 588 1835
rect 535 1767 546 1801
rect 580 1767 588 1801
rect 535 1733 588 1767
rect 535 1699 546 1733
rect 580 1699 588 1733
rect 535 1665 588 1699
rect 535 1631 546 1665
rect 580 1631 588 1665
rect 535 1597 588 1631
rect 535 1563 546 1597
rect 580 1563 588 1597
rect 535 1529 588 1563
rect 535 1495 546 1529
rect 580 1495 588 1529
rect 535 1483 588 1495
rect 362 1292 415 1362
rect 362 1258 370 1292
rect 404 1258 415 1292
rect 362 1224 415 1258
rect 362 1190 370 1224
rect 404 1190 415 1224
rect 362 1156 415 1190
rect 362 1122 370 1156
rect 404 1122 415 1156
rect 362 1088 415 1122
rect 362 1054 370 1088
rect 404 1054 415 1088
rect 362 1020 415 1054
rect 362 986 370 1020
rect 404 986 415 1020
rect 362 952 415 986
rect 362 918 370 952
rect 404 918 415 952
rect 362 884 415 918
rect 362 850 370 884
rect 404 850 415 884
rect 362 816 415 850
rect 362 782 370 816
rect 404 782 415 816
rect 362 748 415 782
rect 362 714 370 748
rect 404 714 415 748
rect 362 680 415 714
rect 362 646 370 680
rect 404 646 415 680
rect 362 612 415 646
rect 362 578 370 612
rect 404 578 415 612
rect 362 544 415 578
rect 362 510 370 544
rect 404 510 415 544
rect 362 476 415 510
rect 362 442 370 476
rect 404 442 415 476
rect 362 408 415 442
rect 362 374 370 408
rect 404 374 415 408
rect 362 362 415 374
rect 535 1292 588 1362
rect 535 1258 546 1292
rect 580 1258 588 1292
rect 535 1224 588 1258
rect 535 1190 546 1224
rect 580 1190 588 1224
rect 535 1156 588 1190
rect 535 1122 546 1156
rect 580 1122 588 1156
rect 535 1088 588 1122
rect 535 1054 546 1088
rect 580 1054 588 1088
rect 535 1020 588 1054
rect 535 986 546 1020
rect 580 986 588 1020
rect 535 952 588 986
rect 535 918 546 952
rect 580 918 588 952
rect 535 884 588 918
rect 535 850 546 884
rect 580 850 588 884
rect 535 816 588 850
rect 535 782 546 816
rect 580 782 588 816
rect 535 748 588 782
rect 535 714 546 748
rect 580 714 588 748
rect 535 680 588 714
rect 535 646 546 680
rect 580 646 588 680
rect 535 612 588 646
rect 535 578 546 612
rect 580 578 588 612
rect 535 544 588 578
rect 535 510 546 544
rect 580 510 588 544
rect 535 476 588 510
rect 535 442 546 476
rect 580 442 588 476
rect 535 408 588 442
rect 535 374 546 408
rect 580 374 588 408
rect 535 362 588 374
<< mvndiffc >>
rect 370 6910 404 6944
rect 370 6842 404 6876
rect 370 6774 404 6808
rect 370 6706 404 6740
rect 370 6638 404 6672
rect 370 6570 404 6604
rect 370 6502 404 6536
rect 370 6434 404 6468
rect 370 6366 404 6400
rect 370 6298 404 6332
rect 370 6230 404 6264
rect 370 6162 404 6196
rect 370 6094 404 6128
rect 370 6026 404 6060
rect 546 6910 580 6944
rect 546 6842 580 6876
rect 546 6774 580 6808
rect 546 6706 580 6740
rect 546 6638 580 6672
rect 546 6570 580 6604
rect 546 6502 580 6536
rect 546 6434 580 6468
rect 546 6366 580 6400
rect 546 6298 580 6332
rect 546 6230 580 6264
rect 546 6162 580 6196
rect 546 6094 580 6128
rect 546 6026 580 6060
rect 370 5789 404 5823
rect 370 5721 404 5755
rect 370 5653 404 5687
rect 370 5585 404 5619
rect 370 5517 404 5551
rect 370 5449 404 5483
rect 370 5381 404 5415
rect 370 5313 404 5347
rect 370 5245 404 5279
rect 370 5177 404 5211
rect 370 5109 404 5143
rect 370 5041 404 5075
rect 370 4973 404 5007
rect 370 4905 404 4939
rect 546 5789 580 5823
rect 546 5721 580 5755
rect 546 5653 580 5687
rect 546 5585 580 5619
rect 546 5517 580 5551
rect 546 5449 580 5483
rect 546 5381 580 5415
rect 546 5313 580 5347
rect 546 5245 580 5279
rect 546 5177 580 5211
rect 546 5109 580 5143
rect 546 5041 580 5075
rect 546 4973 580 5007
rect 546 4905 580 4939
rect 370 4668 404 4702
rect 370 4600 404 4634
rect 370 4532 404 4566
rect 370 4464 404 4498
rect 370 4396 404 4430
rect 370 4328 404 4362
rect 370 4260 404 4294
rect 370 4192 404 4226
rect 370 4124 404 4158
rect 370 4056 404 4090
rect 370 3988 404 4022
rect 370 3920 404 3954
rect 370 3852 404 3886
rect 370 3784 404 3818
rect 546 4668 580 4702
rect 546 4600 580 4634
rect 546 4532 580 4566
rect 546 4464 580 4498
rect 546 4396 580 4430
rect 546 4328 580 4362
rect 546 4260 580 4294
rect 546 4192 580 4226
rect 546 4124 580 4158
rect 546 4056 580 4090
rect 546 3988 580 4022
rect 546 3920 580 3954
rect 546 3852 580 3886
rect 546 3784 580 3818
rect 370 3500 404 3534
rect 370 3432 404 3466
rect 370 3364 404 3398
rect 370 3296 404 3330
rect 370 3228 404 3262
rect 370 3160 404 3194
rect 370 3092 404 3126
rect 370 3024 404 3058
rect 370 2956 404 2990
rect 370 2888 404 2922
rect 370 2820 404 2854
rect 370 2752 404 2786
rect 370 2684 404 2718
rect 370 2616 404 2650
rect 546 3500 580 3534
rect 546 3432 580 3466
rect 546 3364 580 3398
rect 546 3296 580 3330
rect 546 3228 580 3262
rect 546 3160 580 3194
rect 546 3092 580 3126
rect 546 3024 580 3058
rect 546 2956 580 2990
rect 546 2888 580 2922
rect 546 2820 580 2854
rect 546 2752 580 2786
rect 546 2684 580 2718
rect 546 2616 580 2650
rect 370 2379 404 2413
rect 370 2311 404 2345
rect 370 2243 404 2277
rect 370 2175 404 2209
rect 370 2107 404 2141
rect 370 2039 404 2073
rect 370 1971 404 2005
rect 370 1903 404 1937
rect 370 1835 404 1869
rect 370 1767 404 1801
rect 370 1699 404 1733
rect 370 1631 404 1665
rect 370 1563 404 1597
rect 370 1495 404 1529
rect 546 2379 580 2413
rect 546 2311 580 2345
rect 546 2243 580 2277
rect 546 2175 580 2209
rect 546 2107 580 2141
rect 546 2039 580 2073
rect 546 1971 580 2005
rect 546 1903 580 1937
rect 546 1835 580 1869
rect 546 1767 580 1801
rect 546 1699 580 1733
rect 546 1631 580 1665
rect 546 1563 580 1597
rect 546 1495 580 1529
rect 370 1258 404 1292
rect 370 1190 404 1224
rect 370 1122 404 1156
rect 370 1054 404 1088
rect 370 986 404 1020
rect 370 918 404 952
rect 370 850 404 884
rect 370 782 404 816
rect 370 714 404 748
rect 370 646 404 680
rect 370 578 404 612
rect 370 510 404 544
rect 370 442 404 476
rect 370 374 404 408
rect 546 1258 580 1292
rect 546 1190 580 1224
rect 546 1122 580 1156
rect 546 1054 580 1088
rect 546 986 580 1020
rect 546 918 580 952
rect 546 850 580 884
rect 546 782 580 816
rect 546 714 580 748
rect 546 646 580 680
rect 546 578 580 612
rect 546 510 580 544
rect 546 442 580 476
rect 546 374 580 408
<< mvpsubdiff >>
rect 254 7030 278 7064
rect 312 7030 391 7064
rect 425 7030 525 7064
rect 559 7040 696 7064
rect 559 7030 662 7040
rect 254 6972 288 7030
rect 662 6971 696 7006
rect 254 6904 288 6938
rect 254 6836 288 6870
rect 254 6768 288 6802
rect 254 6700 288 6734
rect 254 6632 288 6666
rect 254 6564 288 6598
rect 254 6496 288 6530
rect 254 6428 288 6462
rect 254 6360 288 6394
rect 254 6292 288 6326
rect 254 6224 288 6258
rect 254 6156 288 6190
rect 254 6088 288 6122
rect 254 6020 288 6054
rect 254 5952 288 5986
rect 662 6902 696 6937
rect 662 6833 696 6868
rect 662 6764 696 6799
rect 662 6695 696 6730
rect 662 6626 696 6661
rect 662 6557 696 6592
rect 662 6488 696 6523
rect 662 6419 696 6454
rect 662 6350 696 6385
rect 662 6281 696 6316
rect 662 6212 696 6247
rect 662 6143 696 6178
rect 662 6074 696 6109
rect 662 6005 696 6040
rect 254 5884 288 5918
rect 254 5816 288 5850
rect 662 5936 696 5971
rect 662 5867 696 5902
rect 254 5748 288 5782
rect 254 5680 288 5714
rect 254 5612 288 5646
rect 254 5544 288 5578
rect 254 5476 288 5510
rect 254 5408 288 5442
rect 254 5340 288 5374
rect 254 5272 288 5306
rect 254 5204 288 5238
rect 254 5136 288 5170
rect 254 5068 288 5102
rect 254 5000 288 5034
rect 254 4932 288 4966
rect 254 4864 288 4898
rect 662 5798 696 5833
rect 662 5729 696 5764
rect 662 5660 696 5695
rect 662 5591 696 5626
rect 662 5522 696 5557
rect 662 5453 696 5488
rect 662 5384 696 5419
rect 662 5315 696 5350
rect 662 5246 696 5281
rect 662 5177 696 5212
rect 662 5108 696 5143
rect 662 5039 696 5074
rect 662 4970 696 5005
rect 662 4901 696 4936
rect 254 4796 288 4830
rect 254 4728 288 4762
rect 662 4832 696 4867
rect 662 4763 696 4798
rect 254 4659 288 4694
rect 254 4590 288 4625
rect 254 4521 288 4556
rect 254 4452 288 4487
rect 254 4383 288 4418
rect 254 4314 288 4349
rect 254 4245 288 4280
rect 254 4176 288 4211
rect 254 4107 288 4142
rect 254 4038 288 4073
rect 254 3969 288 4004
rect 254 3900 288 3935
rect 254 3831 288 3866
rect 254 3762 288 3797
rect 254 3693 288 3728
rect 662 4694 696 4729
rect 662 4625 696 4660
rect 662 4556 696 4591
rect 662 4487 696 4522
rect 662 4418 696 4453
rect 662 4349 696 4384
rect 662 4280 696 4315
rect 662 4211 696 4246
rect 662 4142 696 4177
rect 662 4073 696 4108
rect 662 4004 696 4039
rect 662 3935 696 3970
rect 662 3866 696 3901
rect 662 3797 696 3832
rect 662 3728 696 3763
rect 254 3624 288 3659
rect 662 3659 696 3694
rect 254 3555 288 3590
rect 254 3486 288 3521
rect 254 3417 288 3452
rect 254 3348 288 3383
rect 254 3279 288 3314
rect 254 3210 288 3245
rect 254 3141 288 3176
rect 254 3072 288 3107
rect 254 3003 288 3038
rect 254 2934 288 2969
rect 254 2865 288 2900
rect 254 2796 288 2831
rect 254 2727 288 2762
rect 254 2658 288 2693
rect 254 2589 288 2624
rect 662 3590 696 3625
rect 662 3521 696 3556
rect 662 3452 696 3487
rect 662 3383 696 3418
rect 662 3314 696 3349
rect 662 3245 696 3280
rect 662 3176 696 3211
rect 662 3107 696 3142
rect 662 3038 696 3073
rect 662 2969 696 3004
rect 662 2900 696 2935
rect 662 2831 696 2866
rect 662 2762 696 2797
rect 662 2693 696 2728
rect 662 2624 696 2659
rect 254 2520 288 2555
rect 254 2451 288 2486
rect 662 2556 696 2590
rect 662 2488 696 2522
rect 254 2382 288 2417
rect 254 2313 288 2348
rect 254 2244 288 2279
rect 254 2175 288 2210
rect 254 2106 288 2141
rect 254 2037 288 2072
rect 254 1968 288 2003
rect 254 1899 288 1934
rect 254 1830 288 1865
rect 254 1761 288 1796
rect 254 1692 288 1727
rect 254 1623 288 1658
rect 254 1554 288 1589
rect 254 1485 288 1520
rect 662 2420 696 2454
rect 662 2352 696 2386
rect 662 2284 696 2318
rect 662 2216 696 2250
rect 662 2148 696 2182
rect 662 2080 696 2114
rect 662 2012 696 2046
rect 662 1944 696 1978
rect 662 1876 696 1910
rect 662 1808 696 1842
rect 662 1740 696 1774
rect 662 1672 696 1706
rect 662 1604 696 1638
rect 662 1536 696 1570
rect 254 1416 288 1451
rect 254 1347 288 1382
rect 662 1468 696 1502
rect 662 1400 696 1434
rect 254 1278 288 1313
rect 254 1209 288 1244
rect 254 1140 288 1175
rect 254 1071 288 1106
rect 254 1002 288 1037
rect 254 933 288 968
rect 254 864 288 899
rect 254 795 288 830
rect 254 726 288 761
rect 254 657 288 692
rect 254 588 288 623
rect 254 519 288 554
rect 254 450 288 485
rect 254 381 288 416
rect 662 1332 696 1366
rect 662 1264 696 1298
rect 662 1196 696 1230
rect 662 1128 696 1162
rect 662 1060 696 1094
rect 662 992 696 1026
rect 662 924 696 958
rect 662 856 696 890
rect 662 788 696 822
rect 662 720 696 754
rect 662 652 696 686
rect 662 584 696 618
rect 662 516 696 550
rect 662 448 696 482
rect 662 380 696 414
rect 254 312 288 347
rect 662 288 696 346
rect 288 278 352 288
rect 254 254 352 278
rect 386 254 423 288
rect 457 254 494 288
rect 528 254 566 288
rect 600 254 638 288
rect 672 254 696 288
<< mvnsubdiff >>
rect 68 7217 185 7251
rect 219 7217 261 7251
rect 295 7217 337 7251
rect 371 7217 413 7251
rect 447 7217 488 7251
rect 522 7217 563 7251
rect 597 7217 638 7251
rect 672 7217 713 7251
rect 747 7217 882 7251
rect 68 7101 102 7217
rect 68 7033 102 7067
rect 68 6965 102 6999
rect 68 6897 102 6931
rect 68 6829 102 6863
rect 68 6761 102 6795
rect 68 6693 102 6727
rect 68 6625 102 6659
rect 68 6557 102 6591
rect 68 6489 102 6523
rect 68 6421 102 6455
rect 68 6353 102 6387
rect 68 6285 102 6319
rect 68 6217 102 6251
rect 68 6149 102 6183
rect 68 6081 102 6115
rect 68 6013 102 6047
rect 68 5945 102 5979
rect 68 5877 102 5911
rect 68 5809 102 5843
rect 68 5741 102 5775
rect 68 5673 102 5707
rect 68 5605 102 5639
rect 68 5537 102 5571
rect 68 5469 102 5503
rect 68 5401 102 5435
rect 68 5333 102 5367
rect 68 5265 102 5299
rect 68 5197 102 5231
rect 68 5129 102 5163
rect 68 5061 102 5095
rect 68 4993 102 5027
rect 68 4925 102 4959
rect 68 4857 102 4891
rect 68 4789 102 4823
rect 68 4721 102 4755
rect 68 4653 102 4687
rect 68 4585 102 4619
rect 68 4517 102 4551
rect 68 4449 102 4483
rect 68 4381 102 4415
rect 68 4313 102 4347
rect 68 4245 102 4279
rect 68 4177 102 4211
rect 68 4109 102 4143
rect 68 4041 102 4075
rect 68 3973 102 4007
rect 68 3905 102 3939
rect 68 3837 102 3871
rect 68 3769 102 3803
rect 68 3701 102 3735
rect 68 3633 102 3667
rect 68 3565 102 3599
rect 68 3497 102 3531
rect 68 3429 102 3463
rect 68 3361 102 3395
rect 68 3293 102 3327
rect 68 3225 102 3259
rect 68 3157 102 3191
rect 68 3089 102 3123
rect 68 3021 102 3055
rect 68 2953 102 2987
rect 68 2885 102 2919
rect 68 2817 102 2851
rect 68 2749 102 2783
rect 68 2681 102 2715
rect 68 2613 102 2647
rect 68 2545 102 2579
rect 68 2477 102 2511
rect 68 2409 102 2443
rect 68 2341 102 2375
rect 68 2273 102 2307
rect 68 2205 102 2239
rect 68 2137 102 2171
rect 68 2069 102 2103
rect 68 2001 102 2035
rect 68 1933 102 1967
rect 68 1865 102 1899
rect 68 1797 102 1831
rect 68 1729 102 1763
rect 68 1661 102 1695
rect 68 1593 102 1627
rect 68 1525 102 1559
rect 68 1457 102 1491
rect 68 1389 102 1423
rect 68 1321 102 1355
rect 68 1253 102 1287
rect 68 1185 102 1219
rect 68 1117 102 1151
rect 68 1049 102 1083
rect 68 981 102 1015
rect 68 913 102 947
rect 68 845 102 879
rect 68 777 102 811
rect 68 709 102 743
rect 68 641 102 675
rect 68 573 102 607
rect 68 505 102 539
rect 68 437 102 471
rect 68 369 102 403
rect 68 300 102 335
rect 68 231 102 266
rect 68 24 102 197
rect 179 24 203 41
rect 68 7 203 24
rect 237 7 273 41
rect 307 7 344 41
rect 378 7 415 41
rect 449 7 486 41
rect 520 7 557 41
rect 591 7 628 41
rect 662 7 699 41
rect 733 7 770 41
rect 804 24 828 41
rect 848 24 882 7217
rect 804 7 882 24
rect 68 -10 882 7
<< mvpsubdiffcont >>
rect 278 7030 312 7064
rect 391 7030 425 7064
rect 525 7030 559 7064
rect 662 7006 696 7040
rect 254 6938 288 6972
rect 254 6870 288 6904
rect 254 6802 288 6836
rect 254 6734 288 6768
rect 254 6666 288 6700
rect 254 6598 288 6632
rect 254 6530 288 6564
rect 254 6462 288 6496
rect 254 6394 288 6428
rect 254 6326 288 6360
rect 254 6258 288 6292
rect 254 6190 288 6224
rect 254 6122 288 6156
rect 254 6054 288 6088
rect 254 5986 288 6020
rect 662 6937 696 6971
rect 662 6868 696 6902
rect 662 6799 696 6833
rect 662 6730 696 6764
rect 662 6661 696 6695
rect 662 6592 696 6626
rect 662 6523 696 6557
rect 662 6454 696 6488
rect 662 6385 696 6419
rect 662 6316 696 6350
rect 662 6247 696 6281
rect 662 6178 696 6212
rect 662 6109 696 6143
rect 662 6040 696 6074
rect 662 5971 696 6005
rect 254 5918 288 5952
rect 254 5850 288 5884
rect 662 5902 696 5936
rect 254 5782 288 5816
rect 254 5714 288 5748
rect 254 5646 288 5680
rect 254 5578 288 5612
rect 254 5510 288 5544
rect 254 5442 288 5476
rect 254 5374 288 5408
rect 254 5306 288 5340
rect 254 5238 288 5272
rect 254 5170 288 5204
rect 254 5102 288 5136
rect 254 5034 288 5068
rect 254 4966 288 5000
rect 254 4898 288 4932
rect 254 4830 288 4864
rect 662 5833 696 5867
rect 662 5764 696 5798
rect 662 5695 696 5729
rect 662 5626 696 5660
rect 662 5557 696 5591
rect 662 5488 696 5522
rect 662 5419 696 5453
rect 662 5350 696 5384
rect 662 5281 696 5315
rect 662 5212 696 5246
rect 662 5143 696 5177
rect 662 5074 696 5108
rect 662 5005 696 5039
rect 662 4936 696 4970
rect 662 4867 696 4901
rect 254 4762 288 4796
rect 254 4694 288 4728
rect 662 4798 696 4832
rect 662 4729 696 4763
rect 254 4625 288 4659
rect 254 4556 288 4590
rect 254 4487 288 4521
rect 254 4418 288 4452
rect 254 4349 288 4383
rect 254 4280 288 4314
rect 254 4211 288 4245
rect 254 4142 288 4176
rect 254 4073 288 4107
rect 254 4004 288 4038
rect 254 3935 288 3969
rect 254 3866 288 3900
rect 254 3797 288 3831
rect 254 3728 288 3762
rect 662 4660 696 4694
rect 662 4591 696 4625
rect 662 4522 696 4556
rect 662 4453 696 4487
rect 662 4384 696 4418
rect 662 4315 696 4349
rect 662 4246 696 4280
rect 662 4177 696 4211
rect 662 4108 696 4142
rect 662 4039 696 4073
rect 662 3970 696 4004
rect 662 3901 696 3935
rect 662 3832 696 3866
rect 662 3763 696 3797
rect 254 3659 288 3693
rect 254 3590 288 3624
rect 662 3694 696 3728
rect 662 3625 696 3659
rect 254 3521 288 3555
rect 254 3452 288 3486
rect 254 3383 288 3417
rect 254 3314 288 3348
rect 254 3245 288 3279
rect 254 3176 288 3210
rect 254 3107 288 3141
rect 254 3038 288 3072
rect 254 2969 288 3003
rect 254 2900 288 2934
rect 254 2831 288 2865
rect 254 2762 288 2796
rect 254 2693 288 2727
rect 254 2624 288 2658
rect 662 3556 696 3590
rect 662 3487 696 3521
rect 662 3418 696 3452
rect 662 3349 696 3383
rect 662 3280 696 3314
rect 662 3211 696 3245
rect 662 3142 696 3176
rect 662 3073 696 3107
rect 662 3004 696 3038
rect 662 2935 696 2969
rect 662 2866 696 2900
rect 662 2797 696 2831
rect 662 2728 696 2762
rect 662 2659 696 2693
rect 254 2555 288 2589
rect 254 2486 288 2520
rect 662 2590 696 2624
rect 662 2522 696 2556
rect 254 2417 288 2451
rect 254 2348 288 2382
rect 254 2279 288 2313
rect 254 2210 288 2244
rect 254 2141 288 2175
rect 254 2072 288 2106
rect 254 2003 288 2037
rect 254 1934 288 1968
rect 254 1865 288 1899
rect 254 1796 288 1830
rect 254 1727 288 1761
rect 254 1658 288 1692
rect 254 1589 288 1623
rect 254 1520 288 1554
rect 254 1451 288 1485
rect 662 2454 696 2488
rect 662 2386 696 2420
rect 662 2318 696 2352
rect 662 2250 696 2284
rect 662 2182 696 2216
rect 662 2114 696 2148
rect 662 2046 696 2080
rect 662 1978 696 2012
rect 662 1910 696 1944
rect 662 1842 696 1876
rect 662 1774 696 1808
rect 662 1706 696 1740
rect 662 1638 696 1672
rect 662 1570 696 1604
rect 662 1502 696 1536
rect 254 1382 288 1416
rect 662 1434 696 1468
rect 662 1366 696 1400
rect 254 1313 288 1347
rect 254 1244 288 1278
rect 254 1175 288 1209
rect 254 1106 288 1140
rect 254 1037 288 1071
rect 254 968 288 1002
rect 254 899 288 933
rect 254 830 288 864
rect 254 761 288 795
rect 254 692 288 726
rect 254 623 288 657
rect 254 554 288 588
rect 254 485 288 519
rect 254 416 288 450
rect 254 347 288 381
rect 662 1298 696 1332
rect 662 1230 696 1264
rect 662 1162 696 1196
rect 662 1094 696 1128
rect 662 1026 696 1060
rect 662 958 696 992
rect 662 890 696 924
rect 662 822 696 856
rect 662 754 696 788
rect 662 686 696 720
rect 662 618 696 652
rect 662 550 696 584
rect 662 482 696 516
rect 662 414 696 448
rect 662 346 696 380
rect 254 278 288 312
rect 352 254 386 288
rect 423 254 457 288
rect 494 254 528 288
rect 566 254 600 288
rect 638 254 672 288
<< mvnsubdiffcont >>
rect 185 7217 219 7251
rect 261 7217 295 7251
rect 337 7217 371 7251
rect 413 7217 447 7251
rect 488 7217 522 7251
rect 563 7217 597 7251
rect 638 7217 672 7251
rect 713 7217 747 7251
rect 68 7067 102 7101
rect 68 6999 102 7033
rect 68 6931 102 6965
rect 68 6863 102 6897
rect 68 6795 102 6829
rect 68 6727 102 6761
rect 68 6659 102 6693
rect 68 6591 102 6625
rect 68 6523 102 6557
rect 68 6455 102 6489
rect 68 6387 102 6421
rect 68 6319 102 6353
rect 68 6251 102 6285
rect 68 6183 102 6217
rect 68 6115 102 6149
rect 68 6047 102 6081
rect 68 5979 102 6013
rect 68 5911 102 5945
rect 68 5843 102 5877
rect 68 5775 102 5809
rect 68 5707 102 5741
rect 68 5639 102 5673
rect 68 5571 102 5605
rect 68 5503 102 5537
rect 68 5435 102 5469
rect 68 5367 102 5401
rect 68 5299 102 5333
rect 68 5231 102 5265
rect 68 5163 102 5197
rect 68 5095 102 5129
rect 68 5027 102 5061
rect 68 4959 102 4993
rect 68 4891 102 4925
rect 68 4823 102 4857
rect 68 4755 102 4789
rect 68 4687 102 4721
rect 68 4619 102 4653
rect 68 4551 102 4585
rect 68 4483 102 4517
rect 68 4415 102 4449
rect 68 4347 102 4381
rect 68 4279 102 4313
rect 68 4211 102 4245
rect 68 4143 102 4177
rect 68 4075 102 4109
rect 68 4007 102 4041
rect 68 3939 102 3973
rect 68 3871 102 3905
rect 68 3803 102 3837
rect 68 3735 102 3769
rect 68 3667 102 3701
rect 68 3599 102 3633
rect 68 3531 102 3565
rect 68 3463 102 3497
rect 68 3395 102 3429
rect 68 3327 102 3361
rect 68 3259 102 3293
rect 68 3191 102 3225
rect 68 3123 102 3157
rect 68 3055 102 3089
rect 68 2987 102 3021
rect 68 2919 102 2953
rect 68 2851 102 2885
rect 68 2783 102 2817
rect 68 2715 102 2749
rect 68 2647 102 2681
rect 68 2579 102 2613
rect 68 2511 102 2545
rect 68 2443 102 2477
rect 68 2375 102 2409
rect 68 2307 102 2341
rect 68 2239 102 2273
rect 68 2171 102 2205
rect 68 2103 102 2137
rect 68 2035 102 2069
rect 68 1967 102 2001
rect 68 1899 102 1933
rect 68 1831 102 1865
rect 68 1763 102 1797
rect 68 1695 102 1729
rect 68 1627 102 1661
rect 68 1559 102 1593
rect 68 1491 102 1525
rect 68 1423 102 1457
rect 68 1355 102 1389
rect 68 1287 102 1321
rect 68 1219 102 1253
rect 68 1151 102 1185
rect 68 1083 102 1117
rect 68 1015 102 1049
rect 68 947 102 981
rect 68 879 102 913
rect 68 811 102 845
rect 68 743 102 777
rect 68 675 102 709
rect 68 607 102 641
rect 68 539 102 573
rect 68 471 102 505
rect 68 403 102 437
rect 68 335 102 369
rect 68 266 102 300
rect 68 197 102 231
rect 203 7 237 41
rect 273 7 307 41
rect 344 7 378 41
rect 415 7 449 41
rect 486 7 520 41
rect 557 7 591 41
rect 628 7 662 41
rect 699 7 733 41
rect 770 7 804 41
<< poly >>
rect 415 6956 535 6982
rect 415 5916 535 5956
rect 415 5882 472 5916
rect 506 5882 535 5916
rect 415 5835 535 5882
rect 415 4795 535 4835
rect 415 4761 472 4795
rect 506 4761 535 4795
rect 415 4714 535 4761
rect 415 3676 535 3714
rect 415 3642 472 3676
rect 506 3642 535 3676
rect 415 3604 535 3642
rect 415 2556 535 2604
rect 415 2522 472 2556
rect 506 2522 535 2556
rect 415 2483 535 2522
rect 415 1435 535 1483
rect 415 1401 472 1435
rect 506 1401 535 1435
rect 415 1362 535 1401
rect 415 336 535 362
<< polycont >>
rect 472 5882 506 5916
rect 472 4761 506 4795
rect 472 3642 506 3676
rect 472 2522 506 2556
rect 472 1401 506 1435
<< locali >>
rect -44 7217 185 7251
rect 219 7217 261 7251
rect 295 7217 337 7251
rect 371 7217 413 7251
rect 447 7217 488 7251
rect 522 7217 563 7251
rect 597 7217 638 7251
rect 672 7217 713 7251
rect 747 7217 882 7251
rect -44 7101 102 7217
rect -44 7067 68 7101
rect -44 7033 102 7067
rect -44 6999 68 7033
rect -44 6965 102 6999
rect -44 6931 68 6965
rect -44 6897 102 6931
rect -44 6863 68 6897
rect -44 6829 102 6863
rect -44 6795 68 6829
rect -44 6761 102 6795
rect -44 6727 68 6761
rect -44 6693 102 6727
rect -44 6659 68 6693
rect -44 6625 102 6659
rect -44 6591 68 6625
rect -44 6557 102 6591
rect -44 6523 68 6557
rect -44 6489 102 6523
rect -44 6455 68 6489
rect -44 6421 102 6455
rect -44 6387 68 6421
rect -44 6353 102 6387
rect -44 6319 68 6353
rect -44 6285 102 6319
rect -44 6251 68 6285
rect -44 6217 102 6251
rect -44 6183 68 6217
rect -44 6149 102 6183
rect -44 6115 68 6149
rect -44 6081 102 6115
rect -44 6047 68 6081
rect -44 6013 102 6047
rect -44 5979 68 6013
rect -44 5945 102 5979
rect -44 5911 68 5945
rect -44 5877 102 5911
rect -44 5843 68 5877
rect -44 5809 102 5843
rect -44 5775 68 5809
rect -44 5741 102 5775
rect -44 5707 68 5741
rect -44 5673 102 5707
rect -44 5639 68 5673
rect -44 5605 102 5639
rect -44 5571 68 5605
rect -44 5537 102 5571
rect -44 5503 68 5537
rect -44 5469 102 5503
rect -44 5435 68 5469
rect -44 5401 102 5435
rect -44 5367 68 5401
rect -44 5333 102 5367
rect -44 5299 68 5333
rect -44 5265 102 5299
rect -44 5231 68 5265
rect -44 5197 102 5231
rect -44 5163 68 5197
rect -44 5129 102 5163
rect -44 5095 68 5129
rect -44 5061 102 5095
rect -44 5027 68 5061
rect -44 4993 102 5027
rect -44 4959 68 4993
rect -44 4925 102 4959
rect -44 4891 68 4925
rect -44 4857 102 4891
rect -44 4823 68 4857
rect -44 4789 102 4823
rect -44 4755 68 4789
rect -44 4721 102 4755
rect -44 4687 68 4721
rect -44 4653 102 4687
rect -44 4619 68 4653
rect -44 4585 102 4619
rect -44 4551 68 4585
rect -44 4517 102 4551
rect -44 4483 68 4517
rect -44 4449 102 4483
rect -44 4415 68 4449
rect -44 4381 102 4415
rect -44 4347 68 4381
rect -44 4313 102 4347
rect -44 4279 68 4313
rect -44 4245 102 4279
rect -44 4211 68 4245
rect -44 4177 102 4211
rect -44 4143 68 4177
rect -44 4109 102 4143
rect -44 4075 68 4109
rect -44 4041 102 4075
rect -44 4007 68 4041
rect -44 3973 102 4007
rect -44 3939 68 3973
rect -44 3905 102 3939
rect -44 3871 68 3905
rect -44 3837 102 3871
rect -44 3803 68 3837
rect -44 3769 102 3803
rect -44 3735 68 3769
rect -44 3701 102 3735
rect -44 3667 68 3701
rect -44 3633 102 3667
rect -44 3599 68 3633
rect -44 3565 102 3599
rect -44 3531 68 3565
rect -44 3497 102 3531
rect -44 3463 68 3497
rect -44 3436 102 3463
rect 24 3429 102 3436
rect 24 3395 68 3429
rect 24 3361 102 3395
rect 24 3327 68 3361
rect 24 3293 102 3327
rect 24 3262 68 3293
rect -35 3259 68 3262
rect -35 3225 102 3259
rect -35 3191 68 3225
rect -35 3157 102 3191
rect -35 3123 68 3157
rect -35 3089 102 3123
rect -35 3055 68 3089
rect -35 3021 102 3055
rect -35 2987 68 3021
rect -35 2953 102 2987
rect -35 2919 68 2953
rect -35 2885 102 2919
rect -35 2851 68 2885
rect -35 2817 102 2851
rect -35 2783 68 2817
rect -35 2749 102 2783
rect -35 2715 68 2749
rect -35 2681 102 2715
rect -35 2647 68 2681
rect -35 2613 102 2647
rect -35 2579 68 2613
rect -35 2545 102 2579
rect -35 2511 68 2545
rect -35 2477 102 2511
rect -35 2443 68 2477
rect -35 2409 102 2443
rect -35 2375 68 2409
rect -35 2341 102 2375
rect -35 2307 68 2341
rect -35 2273 102 2307
rect -35 2239 68 2273
rect -35 2205 102 2239
rect -35 2171 68 2205
rect -35 2137 102 2171
rect -35 2103 68 2137
rect -35 2069 102 2103
rect -35 2035 68 2069
rect -35 2001 102 2035
rect -35 1967 68 2001
rect -35 1933 102 1967
rect -35 1899 68 1933
rect -35 1865 102 1899
rect -35 1831 68 1865
rect -35 1797 102 1831
rect -35 1763 68 1797
rect -35 1729 102 1763
rect -35 1695 68 1729
rect -35 1661 102 1695
rect -35 1627 68 1661
rect -35 1593 102 1627
rect -35 1559 68 1593
rect -35 1525 102 1559
rect -35 1491 68 1525
rect -35 1457 102 1491
rect -35 1423 68 1457
rect -35 1389 102 1423
rect -35 1355 68 1389
rect -35 1321 102 1355
rect -35 1287 68 1321
rect -35 1253 102 1287
rect -35 1219 68 1253
rect -35 1185 102 1219
rect -35 1151 68 1185
rect -35 1117 102 1151
rect -35 1083 68 1117
rect -35 1049 102 1083
rect -35 1015 68 1049
rect -35 981 102 1015
rect -35 947 68 981
rect -35 913 102 947
rect -35 879 68 913
rect -35 845 102 879
rect -35 811 68 845
rect -35 777 102 811
rect -35 743 68 777
rect -35 709 102 743
rect -35 675 68 709
rect -35 641 102 675
rect -35 607 68 641
rect -35 573 102 607
rect -35 539 68 573
rect -35 505 102 539
rect -35 471 68 505
rect -35 437 102 471
rect -35 403 68 437
rect -35 369 102 403
rect -35 335 68 369
rect -35 300 102 335
rect -35 266 68 300
rect -35 231 102 266
rect -35 197 68 231
rect -35 32 102 197
rect 154 7064 796 7165
rect 154 7030 278 7064
rect 312 7030 391 7064
rect 425 7030 525 7064
rect 559 7040 796 7064
rect 559 7030 662 7040
rect 154 7006 662 7030
rect 696 7006 796 7040
rect 154 7000 796 7006
rect 154 6972 318 7000
rect 154 6938 254 6972
rect 288 6938 318 6972
rect 523 6971 796 7000
rect 154 6904 318 6938
rect 154 6870 254 6904
rect 288 6899 318 6904
rect 154 6865 284 6870
rect 154 6836 318 6865
rect 154 6802 254 6836
rect 288 6820 318 6836
rect 154 6786 284 6802
rect 154 6768 318 6786
rect 154 6734 254 6768
rect 288 6742 318 6768
rect 154 6708 284 6734
rect 154 6700 318 6708
rect 154 6666 254 6700
rect 288 6666 318 6700
rect 154 6664 318 6666
rect 154 6632 284 6664
rect 154 6598 254 6632
rect 288 6598 318 6630
rect 154 6586 318 6598
rect 154 6564 284 6586
rect 154 6530 254 6564
rect 288 6530 318 6552
rect 154 6508 318 6530
rect 154 6496 284 6508
rect 154 6462 254 6496
rect 288 6462 318 6474
rect 154 6430 318 6462
rect 154 6428 284 6430
rect 154 6394 254 6428
rect 288 6394 318 6396
rect 154 6360 318 6394
rect 154 6326 254 6360
rect 288 6352 318 6360
rect 154 6318 284 6326
rect 154 6292 318 6318
rect 154 6258 254 6292
rect 288 6274 318 6292
rect 154 6240 284 6258
rect 154 6224 318 6240
rect 154 6190 254 6224
rect 288 6196 318 6224
rect 154 6162 284 6190
rect 154 6156 318 6162
rect 154 6122 254 6156
rect 288 6122 318 6156
rect 154 6088 318 6122
rect 154 6054 254 6088
rect 288 6054 318 6088
rect 154 6020 318 6054
rect 154 5986 254 6020
rect 288 5986 318 6020
rect 154 5952 318 5986
rect 154 5918 254 5952
rect 288 5918 318 5952
rect 154 5884 318 5918
rect 154 5850 254 5884
rect 288 5850 318 5884
rect 154 5816 318 5850
rect 154 5782 254 5816
rect 288 5782 318 5816
rect 154 5748 318 5782
rect 154 5714 254 5748
rect 288 5714 318 5748
rect 154 5680 318 5714
rect 154 5646 254 5680
rect 288 5646 318 5680
rect 154 5612 318 5646
rect 154 5578 254 5612
rect 288 5578 318 5612
rect 154 5544 318 5578
rect 154 5510 254 5544
rect 288 5510 318 5544
rect 154 5476 318 5510
rect 154 5442 254 5476
rect 288 5442 318 5476
rect 154 5408 318 5442
rect 154 5374 254 5408
rect 288 5374 318 5408
rect 154 5340 318 5374
rect 154 5306 254 5340
rect 288 5306 318 5340
rect 154 5272 318 5306
rect 154 5238 254 5272
rect 288 5238 318 5272
rect 154 5204 318 5238
rect 154 5170 254 5204
rect 288 5170 318 5204
rect 154 5136 318 5170
rect 154 5102 254 5136
rect 288 5102 318 5136
rect 154 5068 318 5102
rect 154 5034 254 5068
rect 288 5034 318 5068
rect 154 5000 318 5034
rect 154 4966 254 5000
rect 288 4966 318 5000
rect 154 4932 318 4966
rect 154 4898 254 4932
rect 288 4898 318 4932
rect 154 4864 318 4898
rect 154 4830 254 4864
rect 288 4830 318 4864
rect 154 4796 318 4830
rect 154 4762 254 4796
rect 288 4762 318 4796
rect 154 4728 318 4762
rect 154 4694 254 4728
rect 288 4694 318 4728
rect 154 4659 318 4694
rect 154 4625 254 4659
rect 288 4625 318 4659
rect 154 4590 318 4625
rect 154 4556 254 4590
rect 288 4556 318 4590
rect 154 4521 318 4556
rect 154 4487 254 4521
rect 288 4487 318 4521
rect 154 4452 318 4487
rect 154 4418 254 4452
rect 288 4418 318 4452
rect 154 4383 318 4418
rect 154 4349 254 4383
rect 288 4349 318 4383
rect 154 4314 318 4349
rect 154 4280 254 4314
rect 288 4280 318 4314
rect 154 4245 318 4280
rect 154 4211 254 4245
rect 288 4211 318 4245
rect 154 4176 318 4211
rect 154 4142 254 4176
rect 288 4142 318 4176
rect 154 4107 318 4142
rect 154 4073 254 4107
rect 288 4073 318 4107
rect 154 4038 318 4073
rect 154 4004 254 4038
rect 288 4004 318 4038
rect 154 3969 318 4004
rect 154 3935 254 3969
rect 288 3935 318 3969
rect 154 3900 318 3935
rect 154 3866 254 3900
rect 288 3866 318 3900
rect 154 3831 318 3866
rect 154 3797 254 3831
rect 288 3797 318 3831
rect 154 3762 318 3797
rect 154 3728 254 3762
rect 288 3728 318 3762
rect 154 3693 318 3728
rect 154 3659 254 3693
rect 288 3659 318 3693
rect 154 3624 318 3659
rect 154 3590 254 3624
rect 288 3590 318 3624
rect 154 3555 318 3590
rect 154 3521 254 3555
rect 288 3521 318 3555
rect 154 3486 318 3521
rect 154 3452 254 3486
rect 288 3452 318 3486
rect 154 3417 318 3452
rect 154 3383 254 3417
rect 288 3383 318 3417
rect 154 3348 318 3383
rect 154 3314 254 3348
rect 288 3314 318 3348
rect 154 3279 318 3314
rect 154 3245 254 3279
rect 288 3245 318 3279
rect 154 3210 318 3245
rect 154 3176 254 3210
rect 288 3176 318 3210
rect 154 3141 318 3176
rect 154 3107 254 3141
rect 288 3107 318 3141
rect 154 3072 318 3107
rect 154 3038 254 3072
rect 288 3038 318 3072
rect 154 3003 318 3038
rect 154 2969 254 3003
rect 288 2969 318 3003
rect 154 2934 318 2969
rect 154 2900 254 2934
rect 288 2900 318 2934
rect 154 2865 318 2900
rect 154 2831 254 2865
rect 288 2831 318 2865
rect 154 2796 318 2831
rect 154 2762 254 2796
rect 288 2762 318 2796
rect 154 2727 318 2762
rect 154 2693 254 2727
rect 288 2693 318 2727
rect 154 2658 318 2693
rect 154 2624 254 2658
rect 288 2624 318 2658
rect 154 2589 318 2624
rect 154 2555 254 2589
rect 288 2555 318 2589
rect 154 2520 318 2555
rect 154 2486 254 2520
rect 288 2486 318 2520
rect 154 2451 318 2486
rect 154 2417 254 2451
rect 288 2417 318 2451
rect 154 2382 318 2417
rect 154 2348 254 2382
rect 288 2348 318 2382
rect 154 2313 318 2348
rect 154 2279 254 2313
rect 288 2279 318 2313
rect 154 2244 318 2279
rect 154 2210 254 2244
rect 288 2210 318 2244
rect 154 2175 318 2210
rect 154 2141 254 2175
rect 288 2141 318 2175
rect 154 2106 318 2141
rect 154 2072 254 2106
rect 288 2072 318 2106
rect 154 2037 318 2072
rect 154 2003 254 2037
rect 288 2003 318 2037
rect 154 1968 318 2003
rect 154 1934 254 1968
rect 288 1934 318 1968
rect 154 1899 318 1934
rect 154 1865 254 1899
rect 288 1865 318 1899
rect 154 1830 318 1865
rect 154 1796 254 1830
rect 288 1796 318 1830
rect 154 1761 318 1796
rect 154 1727 254 1761
rect 288 1727 318 1761
rect 154 1692 318 1727
rect 154 1658 254 1692
rect 288 1658 318 1692
rect 154 1623 318 1658
rect 154 1589 254 1623
rect 288 1589 318 1623
rect 154 1570 318 1589
rect 154 1554 284 1570
rect 154 1520 254 1554
rect 288 1520 318 1536
rect 154 1496 318 1520
rect 154 1485 284 1496
rect 154 1451 254 1485
rect 288 1451 318 1462
rect 154 1422 318 1451
rect 154 1416 284 1422
rect 154 1382 254 1416
rect 288 1382 318 1388
rect 154 1348 318 1382
rect 154 1347 284 1348
rect 154 1313 254 1347
rect 288 1313 318 1314
rect 154 1278 318 1313
rect 154 1244 254 1278
rect 288 1274 318 1278
rect 154 1240 284 1244
rect 154 1209 318 1240
rect 154 1175 254 1209
rect 288 1200 318 1209
rect 154 1166 284 1175
rect 154 1140 318 1166
rect 154 1106 254 1140
rect 288 1126 318 1140
rect 154 1092 284 1106
rect 154 1071 318 1092
rect 154 1037 254 1071
rect 288 1052 318 1071
rect 154 1018 284 1037
rect 154 1002 318 1018
rect 154 968 254 1002
rect 288 978 318 1002
rect 154 944 284 968
rect 154 933 318 944
rect 154 899 254 933
rect 288 903 318 933
rect 154 869 284 899
rect 154 864 318 869
rect 154 830 254 864
rect 288 830 318 864
rect 154 828 318 830
rect 154 795 284 828
rect 154 761 254 795
rect 288 761 318 794
rect 154 753 318 761
rect 154 726 284 753
rect 154 692 254 726
rect 288 692 318 719
rect 154 678 318 692
rect 154 657 284 678
rect 154 623 254 657
rect 288 623 318 644
rect 154 603 318 623
rect 154 588 284 603
rect 154 554 254 588
rect 288 554 318 569
rect 154 528 318 554
rect 154 519 284 528
rect 154 485 254 519
rect 288 485 318 494
rect 154 453 318 485
rect 154 450 284 453
rect 154 416 254 450
rect 288 416 318 419
rect 154 381 318 416
rect 154 347 254 381
rect 288 347 318 381
rect 370 6944 471 6960
rect 404 6910 471 6944
rect 370 6876 471 6910
rect 404 6842 471 6876
rect 370 6808 471 6842
rect 404 6774 471 6808
rect 370 6740 471 6774
rect 404 6706 471 6740
rect 370 6672 471 6706
rect 404 6638 471 6672
rect 370 6604 471 6638
rect 404 6570 471 6604
rect 370 6536 471 6570
rect 404 6502 471 6536
rect 370 6468 471 6502
rect 404 6434 471 6468
rect 370 6400 471 6434
rect 404 6366 471 6400
rect 370 6332 471 6366
rect 404 6298 471 6332
rect 370 6264 471 6298
rect 404 6230 471 6264
rect 370 6196 471 6230
rect 404 6162 471 6196
rect 370 6128 471 6162
rect 404 6094 471 6128
rect 370 6060 471 6094
rect 404 6026 471 6060
rect 370 5966 471 6026
rect 523 6944 662 6971
rect 523 6910 546 6944
rect 580 6937 662 6944
rect 696 6937 796 6971
rect 580 6910 796 6937
rect 523 6902 796 6910
rect 523 6899 662 6902
rect 523 6842 546 6899
rect 580 6868 662 6899
rect 696 6868 796 6902
rect 580 6842 796 6868
rect 523 6833 796 6842
rect 523 6820 662 6833
rect 523 6774 546 6820
rect 580 6799 662 6820
rect 696 6799 796 6833
rect 580 6774 796 6799
rect 523 6764 796 6774
rect 523 6742 662 6764
rect 523 6706 546 6742
rect 580 6730 662 6742
rect 696 6730 796 6764
rect 580 6706 796 6730
rect 523 6695 796 6706
rect 523 6672 662 6695
rect 523 6630 546 6672
rect 580 6661 662 6672
rect 696 6661 796 6695
rect 580 6630 796 6661
rect 523 6626 796 6630
rect 523 6604 662 6626
rect 523 6552 546 6604
rect 580 6592 662 6604
rect 696 6592 796 6626
rect 580 6557 796 6592
rect 580 6552 662 6557
rect 523 6536 662 6552
rect 523 6474 546 6536
rect 580 6523 662 6536
rect 696 6523 796 6557
rect 580 6488 796 6523
rect 580 6474 662 6488
rect 523 6468 662 6474
rect 523 6434 546 6468
rect 580 6454 662 6468
rect 696 6454 796 6488
rect 580 6434 796 6454
rect 523 6430 796 6434
rect 523 6366 546 6430
rect 580 6419 796 6430
rect 580 6385 662 6419
rect 696 6385 796 6419
rect 580 6366 796 6385
rect 523 6352 796 6366
rect 523 6298 546 6352
rect 580 6350 796 6352
rect 580 6316 662 6350
rect 696 6316 796 6350
rect 580 6298 796 6316
rect 523 6281 796 6298
rect 523 6274 662 6281
rect 523 6230 546 6274
rect 580 6247 662 6274
rect 696 6247 796 6281
rect 580 6230 796 6247
rect 523 6212 796 6230
rect 523 6196 662 6212
rect 523 6162 546 6196
rect 580 6178 662 6196
rect 696 6178 796 6212
rect 580 6162 796 6178
rect 523 6143 796 6162
rect 523 6128 662 6143
rect 523 6094 546 6128
rect 580 6109 662 6128
rect 696 6109 796 6143
rect 580 6094 796 6109
rect 523 6074 796 6094
rect 523 6060 662 6074
rect 523 6026 546 6060
rect 580 6040 662 6060
rect 696 6040 796 6074
rect 580 6026 796 6040
rect 523 6005 796 6026
rect 523 5971 662 6005
rect 696 5971 796 6005
rect 523 5966 796 5971
rect 370 5838 438 5966
rect 546 5936 796 5966
rect 404 5789 438 5838
rect 370 5764 438 5789
rect 404 5721 438 5764
rect 370 5690 438 5721
rect 404 5653 438 5690
rect 370 5619 438 5653
rect 404 5582 438 5619
rect 370 5551 438 5582
rect 404 5508 438 5551
rect 370 5483 438 5508
rect 404 5434 438 5483
rect 370 5415 438 5434
rect 404 5360 438 5415
rect 370 5347 438 5360
rect 404 5285 438 5347
rect 370 5279 438 5285
rect 404 5245 438 5279
rect 370 5244 438 5245
rect 404 5177 438 5244
rect 370 5169 438 5177
rect 404 5109 438 5169
rect 370 5094 438 5109
rect 404 5041 438 5094
rect 370 5019 438 5041
rect 404 4973 438 5019
rect 370 4944 438 4973
rect 404 4905 438 4944
rect 370 4869 438 4905
rect 404 4835 438 4869
rect 370 4794 438 4835
rect 404 4760 438 4794
rect 370 4702 438 4760
rect 404 4668 438 4702
rect 370 4634 438 4668
rect 404 4600 438 4634
rect 370 4566 438 4600
rect 404 4532 438 4566
rect 370 4498 438 4532
rect 404 4464 438 4498
rect 370 4430 438 4464
rect 404 4396 438 4430
rect 370 4362 438 4396
rect 404 4328 438 4362
rect 370 4294 438 4328
rect 404 4260 438 4294
rect 370 4226 438 4260
rect 404 4192 438 4226
rect 370 4158 438 4192
rect 404 4124 438 4158
rect 370 4090 438 4124
rect 404 4056 438 4090
rect 370 4022 438 4056
rect 404 3988 438 4022
rect 370 3954 438 3988
rect 404 3920 438 3954
rect 370 3886 438 3920
rect 404 3852 438 3886
rect 370 3818 438 3852
rect 404 3784 438 3818
rect 370 3534 438 3784
rect 404 3500 438 3534
rect 370 3466 438 3500
rect 404 3432 438 3466
rect 370 3398 438 3432
rect 404 3364 438 3398
rect 370 3330 438 3364
rect 404 3296 438 3330
rect 370 3262 438 3296
rect 404 3228 438 3262
rect 370 3194 438 3228
rect 404 3160 438 3194
rect 370 3126 438 3160
rect 404 3092 438 3126
rect 370 3058 438 3092
rect 404 3024 438 3058
rect 370 2990 438 3024
rect 404 2938 438 2990
rect 370 2922 438 2938
rect 404 2863 438 2922
rect 370 2854 438 2863
rect 404 2788 438 2854
rect 370 2786 438 2788
rect 404 2752 438 2786
rect 370 2747 438 2752
rect 404 2684 438 2747
rect 370 2672 438 2684
rect 404 2616 438 2672
rect 370 2597 438 2616
rect 404 2563 438 2597
rect 370 2522 438 2563
rect 404 2488 438 2522
rect 370 2447 438 2488
rect 404 2379 438 2447
rect 370 2372 438 2379
rect 404 2311 438 2372
rect 370 2298 438 2311
rect 404 2243 438 2298
rect 370 2224 438 2243
rect 404 2175 438 2224
rect 370 2150 438 2175
rect 404 2107 438 2150
rect 370 2076 438 2107
rect 404 2039 438 2076
rect 370 2005 438 2039
rect 404 1968 438 2005
rect 370 1937 438 1968
rect 404 1894 438 1937
rect 370 1869 438 1894
rect 404 1835 438 1869
rect 370 1801 438 1835
rect 404 1767 438 1801
rect 370 1733 438 1767
rect 404 1699 438 1733
rect 370 1665 438 1699
rect 404 1631 438 1665
rect 370 1597 438 1631
rect 404 1563 438 1597
rect 370 1529 438 1563
rect 404 1495 438 1529
rect 370 1351 438 1495
rect 472 5916 506 5932
rect 472 4795 506 5882
rect 472 4436 506 4761
rect 472 4364 506 4402
rect 472 3676 506 4330
rect 472 3402 506 3642
rect 472 3330 506 3368
rect 472 2556 506 3296
rect 472 1435 506 2522
rect 472 1385 506 1401
rect 546 5902 662 5936
rect 696 5902 796 5936
rect 546 5867 796 5902
rect 546 5833 662 5867
rect 696 5833 796 5867
rect 546 5823 796 5833
rect 580 5798 796 5823
rect 580 5789 662 5798
rect 546 5764 662 5789
rect 696 5764 796 5798
rect 546 5755 796 5764
rect 580 5729 796 5755
rect 580 5721 662 5729
rect 546 5695 662 5721
rect 696 5695 796 5729
rect 546 5687 796 5695
rect 580 5660 796 5687
rect 580 5653 662 5660
rect 546 5626 662 5653
rect 696 5626 796 5660
rect 546 5619 796 5626
rect 580 5591 796 5619
rect 580 5585 662 5591
rect 546 5557 662 5585
rect 696 5557 796 5591
rect 546 5551 796 5557
rect 580 5522 796 5551
rect 580 5517 662 5522
rect 546 5488 662 5517
rect 696 5488 796 5522
rect 546 5483 796 5488
rect 580 5453 796 5483
rect 580 5449 662 5453
rect 546 5419 662 5449
rect 696 5419 796 5453
rect 546 5415 796 5419
rect 580 5384 796 5415
rect 580 5381 662 5384
rect 546 5350 662 5381
rect 696 5350 796 5384
rect 546 5347 796 5350
rect 580 5315 796 5347
rect 580 5313 662 5315
rect 546 5281 662 5313
rect 696 5281 796 5315
rect 546 5279 796 5281
rect 580 5246 796 5279
rect 580 5245 662 5246
rect 546 5212 662 5245
rect 696 5212 796 5246
rect 546 5211 796 5212
rect 580 5177 796 5211
rect 546 5143 662 5177
rect 696 5143 796 5177
rect 580 5109 796 5143
rect 546 5108 796 5109
rect 546 5075 662 5108
rect 580 5074 662 5075
rect 696 5074 796 5108
rect 580 5041 796 5074
rect 546 5039 796 5041
rect 546 5007 662 5039
rect 580 5005 662 5007
rect 696 5005 796 5039
rect 580 4973 796 5005
rect 546 4970 796 4973
rect 546 4939 662 4970
rect 580 4936 662 4939
rect 696 4936 796 4970
rect 580 4905 796 4936
rect 546 4901 796 4905
rect 546 4867 662 4901
rect 696 4867 796 4901
rect 546 4832 796 4867
rect 546 4798 662 4832
rect 696 4798 796 4832
rect 546 4763 796 4798
rect 546 4729 662 4763
rect 696 4729 796 4763
rect 546 4702 796 4729
rect 580 4694 796 4702
rect 580 4668 662 4694
rect 546 4660 662 4668
rect 696 4660 796 4694
rect 546 4634 796 4660
rect 580 4625 796 4634
rect 580 4600 662 4625
rect 546 4591 662 4600
rect 696 4591 796 4625
rect 546 4566 796 4591
rect 580 4556 796 4566
rect 580 4532 662 4556
rect 546 4522 662 4532
rect 696 4522 796 4556
rect 546 4498 796 4522
rect 580 4487 796 4498
rect 580 4464 662 4487
rect 546 4453 662 4464
rect 696 4453 796 4487
rect 546 4430 796 4453
rect 580 4418 796 4430
rect 580 4396 662 4418
rect 546 4384 662 4396
rect 696 4384 796 4418
rect 546 4362 796 4384
rect 580 4349 796 4362
rect 580 4328 662 4349
rect 546 4315 662 4328
rect 696 4315 796 4349
rect 546 4294 796 4315
rect 580 4280 796 4294
rect 580 4260 662 4280
rect 546 4246 662 4260
rect 696 4246 796 4280
rect 546 4226 796 4246
rect 580 4211 796 4226
rect 580 4192 662 4211
rect 546 4177 662 4192
rect 696 4177 796 4211
rect 546 4158 796 4177
rect 580 4142 796 4158
rect 580 4124 662 4142
rect 546 4108 662 4124
rect 696 4108 796 4142
rect 546 4090 796 4108
rect 580 4073 796 4090
rect 580 4056 662 4073
rect 546 4039 662 4056
rect 696 4039 796 4073
rect 546 4022 796 4039
rect 580 4004 796 4022
rect 580 3972 662 4004
rect 546 3970 662 3972
rect 696 3970 796 4004
rect 546 3954 796 3970
rect 580 3935 796 3954
rect 580 3901 662 3935
rect 696 3901 796 3935
rect 580 3890 796 3901
rect 546 3886 796 3890
rect 580 3866 796 3886
rect 580 3852 662 3866
rect 546 3842 662 3852
rect 580 3832 662 3842
rect 696 3832 796 3866
rect 580 3797 796 3832
rect 580 3784 662 3797
rect 546 3763 662 3784
rect 696 3763 796 3797
rect 546 3760 796 3763
rect 580 3728 796 3760
rect 580 3726 662 3728
rect 546 3694 662 3726
rect 696 3694 796 3728
rect 546 3659 796 3694
rect 546 3625 662 3659
rect 696 3625 796 3659
rect 546 3590 796 3625
rect 546 3556 662 3590
rect 696 3556 796 3590
rect 546 3534 796 3556
rect 580 3521 796 3534
rect 580 3500 662 3521
rect 546 3487 662 3500
rect 696 3487 796 3521
rect 546 3466 796 3487
rect 580 3452 796 3466
rect 580 3432 662 3452
rect 546 3418 662 3432
rect 696 3418 796 3452
rect 546 3398 796 3418
rect 580 3383 796 3398
rect 580 3364 662 3383
rect 546 3349 662 3364
rect 696 3349 796 3383
rect 546 3330 796 3349
rect 580 3314 796 3330
rect 580 3296 662 3314
rect 546 3280 662 3296
rect 696 3280 796 3314
rect 546 3262 796 3280
rect 580 3245 796 3262
rect 580 3228 662 3245
rect 546 3211 662 3228
rect 696 3211 796 3245
rect 546 3194 796 3211
rect 580 3176 796 3194
rect 580 3160 662 3176
rect 546 3142 662 3160
rect 696 3142 796 3176
rect 546 3126 796 3142
rect 580 3107 796 3126
rect 580 3092 662 3107
rect 546 3073 662 3092
rect 696 3073 796 3107
rect 546 3058 796 3073
rect 580 3038 796 3058
rect 580 3024 662 3038
rect 546 3004 662 3024
rect 696 3004 796 3038
rect 546 2990 796 3004
rect 580 2969 796 2990
rect 580 2956 662 2969
rect 546 2935 662 2956
rect 696 2935 796 2969
rect 546 2922 796 2935
rect 580 2900 796 2922
rect 580 2888 662 2900
rect 546 2866 662 2888
rect 696 2866 796 2900
rect 546 2854 796 2866
rect 580 2831 796 2854
rect 580 2820 662 2831
rect 546 2797 662 2820
rect 696 2797 796 2831
rect 546 2786 796 2797
rect 580 2762 796 2786
rect 580 2752 662 2762
rect 546 2728 662 2752
rect 696 2728 796 2762
rect 546 2718 796 2728
rect 580 2693 796 2718
rect 580 2684 662 2693
rect 546 2659 662 2684
rect 696 2659 796 2693
rect 546 2650 796 2659
rect 580 2624 796 2650
rect 580 2616 662 2624
rect 546 2590 662 2616
rect 696 2590 796 2624
rect 546 2556 796 2590
rect 546 2522 662 2556
rect 696 2522 796 2556
rect 546 2488 796 2522
rect 546 2454 662 2488
rect 696 2454 796 2488
rect 546 2420 796 2454
rect 546 2413 662 2420
rect 580 2386 662 2413
rect 696 2386 796 2420
rect 580 2379 796 2386
rect 546 2352 796 2379
rect 546 2345 662 2352
rect 580 2318 662 2345
rect 696 2318 796 2352
rect 580 2311 796 2318
rect 546 2284 796 2311
rect 546 2277 662 2284
rect 580 2250 662 2277
rect 696 2250 796 2284
rect 580 2243 796 2250
rect 546 2216 796 2243
rect 546 2209 662 2216
rect 580 2182 662 2209
rect 696 2182 796 2216
rect 580 2175 796 2182
rect 546 2148 796 2175
rect 546 2141 662 2148
rect 580 2114 662 2141
rect 696 2114 796 2148
rect 580 2107 796 2114
rect 546 2080 796 2107
rect 546 2073 662 2080
rect 580 2046 662 2073
rect 696 2046 796 2080
rect 580 2039 796 2046
rect 546 2012 796 2039
rect 546 2005 662 2012
rect 580 1978 662 2005
rect 696 1978 796 2012
rect 580 1971 796 1978
rect 546 1944 796 1971
rect 546 1937 662 1944
rect 580 1910 662 1937
rect 696 1910 796 1944
rect 580 1903 796 1910
rect 546 1876 796 1903
rect 546 1869 662 1876
rect 580 1842 662 1869
rect 696 1842 796 1876
rect 580 1835 796 1842
rect 546 1808 796 1835
rect 546 1801 662 1808
rect 580 1774 662 1801
rect 696 1774 796 1808
rect 580 1767 796 1774
rect 546 1740 796 1767
rect 546 1733 662 1740
rect 580 1706 662 1733
rect 696 1706 796 1740
rect 580 1699 796 1706
rect 546 1672 796 1699
rect 546 1665 662 1672
rect 580 1638 662 1665
rect 696 1638 796 1672
rect 580 1631 796 1638
rect 546 1604 796 1631
rect 546 1597 662 1604
rect 580 1570 662 1597
rect 696 1570 796 1604
rect 580 1563 796 1570
rect 546 1536 796 1563
rect 546 1529 662 1536
rect 580 1502 662 1529
rect 696 1502 796 1536
rect 580 1495 796 1502
rect 546 1468 796 1495
rect 546 1434 662 1468
rect 696 1434 796 1468
rect 546 1400 796 1434
rect 546 1366 662 1400
rect 696 1366 796 1400
rect 546 1351 796 1366
rect 370 1292 471 1351
rect 404 1258 471 1292
rect 370 1224 471 1258
rect 404 1190 471 1224
rect 370 1156 471 1190
rect 404 1122 471 1156
rect 370 1088 471 1122
rect 404 1054 471 1088
rect 370 1020 471 1054
rect 404 986 471 1020
rect 370 952 471 986
rect 404 918 471 952
rect 370 884 471 918
rect 404 850 471 884
rect 370 816 471 850
rect 404 782 471 816
rect 370 748 471 782
rect 404 714 471 748
rect 370 680 471 714
rect 404 646 471 680
rect 370 612 471 646
rect 404 578 471 612
rect 370 544 471 578
rect 404 510 471 544
rect 370 476 471 510
rect 404 442 471 476
rect 370 408 471 442
rect 404 374 471 408
rect 370 358 471 374
rect 523 1317 546 1351
rect 580 1332 796 1351
rect 580 1317 662 1332
rect 523 1298 662 1317
rect 696 1298 796 1332
rect 523 1292 796 1298
rect 523 1243 546 1292
rect 580 1264 796 1292
rect 580 1243 662 1264
rect 523 1230 662 1243
rect 696 1230 796 1264
rect 523 1224 796 1230
rect 523 1169 546 1224
rect 580 1196 796 1224
rect 580 1169 662 1196
rect 523 1162 662 1169
rect 696 1162 796 1196
rect 523 1156 796 1162
rect 523 1094 546 1156
rect 580 1128 796 1156
rect 580 1094 662 1128
rect 696 1094 796 1128
rect 523 1088 796 1094
rect 523 1054 546 1088
rect 580 1060 796 1088
rect 580 1054 662 1060
rect 523 1053 662 1054
rect 523 986 546 1053
rect 580 1026 662 1053
rect 696 1026 796 1060
rect 580 992 796 1026
rect 580 986 662 992
rect 523 978 662 986
rect 523 918 546 978
rect 580 958 662 978
rect 696 958 796 992
rect 580 924 796 958
rect 580 918 662 924
rect 523 903 662 918
rect 523 850 546 903
rect 580 890 662 903
rect 696 890 796 924
rect 580 856 796 890
rect 580 850 662 856
rect 523 828 662 850
rect 523 782 546 828
rect 580 822 662 828
rect 696 822 796 856
rect 580 788 796 822
rect 580 782 662 788
rect 523 754 662 782
rect 696 754 796 788
rect 523 753 796 754
rect 523 714 546 753
rect 580 720 796 753
rect 580 714 662 720
rect 523 686 662 714
rect 696 686 796 720
rect 523 680 796 686
rect 523 644 546 680
rect 580 652 796 680
rect 580 644 662 652
rect 523 618 662 644
rect 696 618 796 652
rect 523 612 796 618
rect 523 569 546 612
rect 580 584 796 612
rect 580 569 662 584
rect 523 550 662 569
rect 696 550 796 584
rect 523 544 796 550
rect 523 494 546 544
rect 580 516 796 544
rect 580 494 662 516
rect 523 482 662 494
rect 696 482 796 516
rect 523 476 796 482
rect 523 419 546 476
rect 580 448 796 476
rect 580 419 662 448
rect 523 414 662 419
rect 696 414 796 448
rect 523 408 796 414
rect 523 374 546 408
rect 580 380 796 408
rect 580 374 662 380
rect 154 318 318 347
rect 523 346 662 374
rect 696 346 796 380
rect 523 318 796 346
rect 154 312 796 318
rect 154 278 254 312
rect 288 288 796 312
rect 288 278 352 288
rect 154 254 352 278
rect 386 254 423 288
rect 457 254 494 288
rect 528 254 566 288
rect 600 254 638 288
rect 672 254 796 288
rect 154 153 796 254
rect 179 32 203 41
rect 237 32 273 41
rect 307 32 344 41
rect -35 -2 28 32
rect 62 -2 106 32
rect 140 -2 184 32
rect 237 7 262 32
rect 307 7 340 32
rect 378 7 415 41
rect 449 32 486 41
rect 520 32 557 41
rect 591 32 628 41
rect 662 32 699 41
rect 733 32 770 41
rect 452 7 486 32
rect 530 7 557 32
rect 608 7 628 32
rect 686 7 699 32
rect 764 7 770 32
rect 804 32 828 41
rect 804 7 808 32
rect 218 -2 262 7
rect 296 -2 340 7
rect 374 -2 418 7
rect 452 -2 496 7
rect 530 -2 574 7
rect 608 -2 652 7
rect 686 -2 730 7
rect 764 -2 808 7
rect 848 24 882 7217
rect 842 -2 882 24
rect -35 -10 882 -2
<< viali >>
rect 284 6870 288 6899
rect 288 6870 318 6899
rect 284 6865 318 6870
rect 284 6802 288 6820
rect 288 6802 318 6820
rect 284 6786 318 6802
rect 284 6734 288 6742
rect 288 6734 318 6742
rect 284 6708 318 6734
rect 284 6632 318 6664
rect 284 6630 288 6632
rect 288 6630 318 6632
rect 284 6564 318 6586
rect 284 6552 288 6564
rect 288 6552 318 6564
rect 284 6496 318 6508
rect 284 6474 288 6496
rect 288 6474 318 6496
rect 284 6428 318 6430
rect 284 6396 288 6428
rect 288 6396 318 6428
rect 284 6326 288 6352
rect 288 6326 318 6352
rect 284 6318 318 6326
rect 284 6258 288 6274
rect 288 6258 318 6274
rect 284 6240 318 6258
rect 284 6190 288 6196
rect 288 6190 318 6196
rect 284 6162 318 6190
rect 284 1554 318 1570
rect 284 1536 288 1554
rect 288 1536 318 1554
rect 284 1485 318 1496
rect 284 1462 288 1485
rect 288 1462 318 1485
rect 284 1416 318 1422
rect 284 1388 288 1416
rect 288 1388 318 1416
rect 284 1347 318 1348
rect 284 1314 288 1347
rect 288 1314 318 1347
rect 284 1244 288 1274
rect 288 1244 318 1274
rect 284 1240 318 1244
rect 284 1175 288 1200
rect 288 1175 318 1200
rect 284 1166 318 1175
rect 284 1106 288 1126
rect 288 1106 318 1126
rect 284 1092 318 1106
rect 284 1037 288 1052
rect 288 1037 318 1052
rect 284 1018 318 1037
rect 284 968 288 978
rect 288 968 318 978
rect 284 944 318 968
rect 284 899 288 903
rect 288 899 318 903
rect 284 869 318 899
rect 284 795 318 828
rect 284 794 288 795
rect 288 794 318 795
rect 284 726 318 753
rect 284 719 288 726
rect 288 719 318 726
rect 284 657 318 678
rect 284 644 288 657
rect 288 644 318 657
rect 284 588 318 603
rect 284 569 288 588
rect 288 569 318 588
rect 284 519 318 528
rect 284 494 288 519
rect 288 494 318 519
rect 284 450 318 453
rect 284 419 288 450
rect 288 419 318 450
rect 546 6876 580 6899
rect 546 6865 580 6876
rect 546 6808 580 6820
rect 546 6786 580 6808
rect 546 6740 580 6742
rect 546 6708 580 6740
rect 546 6638 580 6664
rect 546 6630 580 6638
rect 546 6570 580 6586
rect 546 6552 580 6570
rect 546 6502 580 6508
rect 546 6474 580 6502
rect 546 6400 580 6430
rect 546 6396 580 6400
rect 546 6332 580 6352
rect 546 6318 580 6332
rect 546 6264 580 6274
rect 546 6240 580 6264
rect 546 6162 580 6196
rect 370 5823 404 5838
rect 370 5804 404 5823
rect 370 5755 404 5764
rect 370 5730 404 5755
rect 370 5687 404 5690
rect 370 5656 404 5687
rect 370 5585 404 5616
rect 370 5582 404 5585
rect 370 5517 404 5542
rect 370 5508 404 5517
rect 370 5449 404 5468
rect 370 5434 404 5449
rect 370 5381 404 5394
rect 370 5360 404 5381
rect 370 5313 404 5319
rect 370 5285 404 5313
rect 370 5211 404 5244
rect 370 5210 404 5211
rect 370 5143 404 5169
rect 370 5135 404 5143
rect 370 5075 404 5094
rect 370 5060 404 5075
rect 370 5007 404 5019
rect 370 4985 404 5007
rect 370 4939 404 4944
rect 370 4910 404 4939
rect 370 4835 404 4869
rect 370 4760 404 4794
rect 370 2956 404 2972
rect 370 2938 404 2956
rect 370 2888 404 2897
rect 370 2863 404 2888
rect 370 2820 404 2822
rect 370 2788 404 2820
rect 370 2718 404 2747
rect 370 2713 404 2718
rect 370 2650 404 2672
rect 370 2638 404 2650
rect 370 2563 404 2597
rect 370 2488 404 2522
rect 370 2413 404 2447
rect 370 2345 404 2372
rect 370 2338 404 2345
rect 370 2277 404 2298
rect 370 2264 404 2277
rect 370 2209 404 2224
rect 370 2190 404 2209
rect 370 2141 404 2150
rect 370 2116 404 2141
rect 370 2073 404 2076
rect 370 2042 404 2073
rect 370 1971 404 2002
rect 370 1968 404 1971
rect 370 1903 404 1928
rect 370 1894 404 1903
rect 472 4402 506 4436
rect 472 4330 506 4364
rect 472 3368 506 3402
rect 472 3296 506 3330
rect 546 3988 580 4006
rect 546 3972 580 3988
rect 546 3920 580 3924
rect 546 3890 580 3920
rect 546 3818 580 3842
rect 546 3808 580 3818
rect 546 3726 580 3760
rect 546 1317 580 1351
rect 546 1258 580 1277
rect 546 1243 580 1258
rect 546 1190 580 1203
rect 546 1169 580 1190
rect 546 1122 580 1128
rect 546 1094 580 1122
rect 546 1020 580 1053
rect 546 1019 580 1020
rect 546 952 580 978
rect 546 944 580 952
rect 546 884 580 903
rect 546 869 580 884
rect 546 816 580 828
rect 546 794 580 816
rect 546 748 580 753
rect 546 719 580 748
rect 546 646 580 678
rect 546 644 580 646
rect 546 578 580 603
rect 546 569 580 578
rect 546 510 580 528
rect 546 494 580 510
rect 546 442 580 453
rect 546 419 580 442
rect 28 -2 62 32
rect 106 -2 140 32
rect 184 7 203 32
rect 203 7 218 32
rect 262 7 273 32
rect 273 7 296 32
rect 340 7 344 32
rect 344 7 374 32
rect 418 7 449 32
rect 449 7 452 32
rect 496 7 520 32
rect 520 7 530 32
rect 574 7 591 32
rect 591 7 608 32
rect 652 7 662 32
rect 662 7 686 32
rect 730 7 733 32
rect 733 7 764 32
rect 184 -2 218 7
rect 262 -2 296 7
rect 340 -2 374 7
rect 418 -2 452 7
rect 496 -2 530 7
rect 574 -2 608 7
rect 652 -2 686 7
rect 730 -2 764 7
rect 808 -2 842 32
<< metal1 >>
tri 825 7257 924 7356 se
rect 16 7211 924 7257
tri 833 7120 924 7211 ne
rect 278 6899 586 6911
rect 278 6865 284 6899
rect 318 6865 546 6899
rect 580 6865 586 6899
rect 278 6820 586 6865
rect 278 6786 284 6820
rect 318 6786 546 6820
rect 580 6786 586 6820
rect 278 6742 586 6786
rect 278 6708 284 6742
rect 318 6708 546 6742
rect 580 6708 586 6742
rect 278 6664 586 6708
rect 278 6630 284 6664
rect 318 6630 546 6664
rect 580 6630 586 6664
rect 278 6586 586 6630
rect 278 6552 284 6586
rect 318 6552 546 6586
rect 580 6552 586 6586
rect 278 6508 586 6552
rect 278 6474 284 6508
rect 318 6474 546 6508
rect 580 6474 586 6508
rect 278 6430 586 6474
rect 278 6396 284 6430
rect 318 6396 546 6430
rect 580 6396 586 6430
rect 278 6352 586 6396
rect 278 6318 284 6352
rect 318 6318 546 6352
rect 580 6318 586 6352
rect 278 6274 586 6318
rect 278 6240 284 6274
rect 318 6240 546 6274
rect 580 6240 586 6274
rect 278 6196 586 6240
rect 278 6162 284 6196
rect 318 6162 546 6196
rect 580 6162 586 6196
rect 278 6150 586 6162
rect 364 5838 410 5850
rect 364 5804 370 5838
rect 404 5804 410 5838
rect 364 5764 410 5804
rect 364 5730 370 5764
rect 404 5730 410 5764
rect 364 5690 410 5730
rect 364 5656 370 5690
rect 404 5656 410 5690
rect 364 5616 410 5656
rect 364 5582 370 5616
rect 404 5582 410 5616
rect 364 5542 410 5582
rect 364 5508 370 5542
rect 404 5508 410 5542
rect 364 5468 410 5508
rect 364 5434 370 5468
rect 404 5434 410 5468
rect 364 5394 410 5434
rect 364 5360 370 5394
rect 404 5360 410 5394
rect 364 5319 410 5360
rect 364 5285 370 5319
rect 404 5285 410 5319
rect 364 5244 410 5285
rect 364 5210 370 5244
rect 404 5210 410 5244
rect 364 5169 410 5210
rect 364 5135 370 5169
rect 404 5135 410 5169
rect 364 5094 410 5135
rect 364 5060 370 5094
rect 404 5060 410 5094
rect 364 5019 410 5060
rect 364 4985 370 5019
rect 404 4985 410 5019
rect 364 4944 410 4985
rect 364 4910 370 4944
rect 404 4910 410 4944
tri 339 4878 364 4903 se
rect 364 4878 410 4910
rect -50 4869 410 4878
rect -50 4835 370 4869
rect 404 4835 410 4869
rect -50 4794 410 4835
rect -50 4760 370 4794
rect 404 4760 410 4794
rect -50 4748 410 4760
rect 361 4436 512 4448
rect 361 4402 472 4436
rect 506 4402 512 4436
rect 361 4364 512 4402
rect 361 4330 472 4364
rect 506 4330 512 4364
rect 361 4318 512 4330
rect 278 4018 318 4122
tri 318 4018 422 4122 sw
rect 278 4006 586 4018
rect 278 3972 546 4006
rect 580 3972 586 4006
rect 278 3924 586 3972
rect 278 3890 546 3924
rect 580 3890 586 3924
rect 278 3842 586 3890
rect 278 3808 546 3842
rect 580 3808 586 3842
rect 278 3760 586 3808
rect 278 3726 546 3760
rect 580 3726 586 3760
rect 278 3714 586 3726
rect 278 3608 318 3714
tri 318 3608 424 3714 nw
rect 362 3402 512 3414
rect 362 3368 472 3402
rect 506 3368 512 3402
rect 362 3330 512 3368
rect 362 3296 472 3330
rect 506 3296 512 3330
rect 362 3284 512 3296
rect -50 2972 410 2984
rect -50 2938 370 2972
rect 404 2938 410 2972
rect -50 2897 410 2938
rect -50 2863 370 2897
rect 404 2863 410 2897
rect -50 2854 410 2863
tri 339 2829 364 2854 ne
rect 364 2822 410 2854
rect 364 2788 370 2822
rect 404 2788 410 2822
rect 364 2747 410 2788
rect 364 2713 370 2747
rect 404 2713 410 2747
rect 364 2672 410 2713
rect 364 2638 370 2672
rect 404 2638 410 2672
rect 364 2597 410 2638
rect 364 2563 370 2597
rect 404 2563 410 2597
rect 364 2522 410 2563
rect 364 2488 370 2522
rect 404 2488 410 2522
rect 364 2447 410 2488
rect 364 2413 370 2447
rect 404 2413 410 2447
rect 364 2372 410 2413
rect 364 2338 370 2372
rect 404 2338 410 2372
rect 364 2298 410 2338
rect 364 2264 370 2298
rect 404 2264 410 2298
rect 364 2224 410 2264
rect 364 2190 370 2224
rect 404 2190 410 2224
rect 364 2150 410 2190
rect 364 2116 370 2150
rect 404 2116 410 2150
rect 364 2076 410 2116
rect 364 2042 370 2076
rect 404 2042 410 2076
rect 364 2002 410 2042
rect 364 1968 370 2002
rect 404 1968 410 2002
rect 364 1928 410 1968
rect 364 1894 370 1928
rect 404 1894 410 1928
rect 364 1882 410 1894
rect 278 1570 545 1582
rect 278 1536 284 1570
rect 318 1536 545 1570
rect 278 1496 545 1536
rect 278 1462 284 1496
rect 318 1462 545 1496
rect 278 1422 545 1462
rect 278 1388 284 1422
rect 318 1388 545 1422
rect 278 1363 545 1388
tri 545 1363 586 1404 sw
rect 278 1351 586 1363
rect 278 1348 546 1351
rect 278 1314 284 1348
rect 318 1317 546 1348
rect 580 1317 586 1351
rect 318 1314 586 1317
rect 278 1277 586 1314
rect 278 1274 546 1277
rect 278 1240 284 1274
rect 318 1243 546 1274
rect 580 1243 586 1277
rect 318 1240 586 1243
rect 278 1203 586 1240
rect 278 1200 546 1203
rect 278 1166 284 1200
rect 318 1169 546 1200
rect 580 1169 586 1203
rect 318 1166 586 1169
rect 278 1128 586 1166
rect 278 1126 546 1128
rect 278 1092 284 1126
rect 318 1094 546 1126
rect 580 1094 586 1128
rect 318 1092 586 1094
rect 278 1053 586 1092
rect 278 1052 546 1053
rect 278 1018 284 1052
rect 318 1019 546 1052
rect 580 1019 586 1053
rect 318 1018 586 1019
rect 278 978 586 1018
rect 278 944 284 978
rect 318 944 546 978
rect 580 944 586 978
rect 278 903 586 944
rect 278 869 284 903
rect 318 869 546 903
rect 580 869 586 903
rect 278 828 586 869
rect 278 794 284 828
rect 318 794 546 828
rect 580 794 586 828
rect 278 753 586 794
rect 278 719 284 753
rect 318 719 546 753
rect 580 719 586 753
rect 278 678 586 719
rect 278 644 284 678
rect 318 644 546 678
rect 580 644 586 678
rect 278 603 586 644
rect 278 569 284 603
rect 318 569 546 603
rect 580 569 586 603
rect 278 528 586 569
rect 278 494 284 528
rect 318 494 546 528
rect 580 494 586 528
rect 278 453 586 494
rect 278 419 284 453
rect 318 419 546 453
rect 580 419 586 453
rect 278 407 586 419
tri 856 86 908 138 se
rect 908 86 936 138
rect -26 38 92 86
tri 92 38 140 86 sw
tri 808 38 856 86 se
rect 856 38 936 86
rect -26 32 936 38
rect -26 -2 28 32
rect 62 -2 106 32
rect 140 -2 184 32
rect 218 -2 262 32
rect 296 -2 340 32
rect 374 -2 418 32
rect 452 -2 496 32
rect 530 -2 574 32
rect 608 -2 652 32
rect 686 -2 730 32
rect 764 -2 808 32
rect 842 -2 936 32
rect -26 -8 936 -2
tri 808 -108 908 -8 ne
rect 908 -108 936 -8
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_0
timestamp 1688980957
transform 1 0 415 0 -1 5835
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_1
timestamp 1688980957
transform 1 0 415 0 -1 6956
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_2
timestamp 1688980957
transform 1 0 415 0 1 1483
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_3
timestamp 1688980957
transform 1 0 415 0 1 362
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_4
timestamp 1688980957
transform 1 0 415 0 -1 4714
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_5
timestamp 1688980957
transform 1 0 415 0 1 2604
box -1 0 121 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1688980957
transform 0 -1 506 1 0 3296
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1688980957
transform 0 -1 506 -1 0 4436
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_0
timestamp 1688980957
transform 1 0 456 0 1 1385
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_1
timestamp 1688980957
transform 1 0 456 0 1 3626
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_2
timestamp 1688980957
transform 1 0 456 0 1 5866
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_3
timestamp 1688980957
transform 1 0 456 0 1 4745
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_4
timestamp 1688980957
transform 1 0 456 0 1 2506
box 0 0 1 1
<< labels >>
flabel comment s 229 6177 229 6177 0 FreeSans 400 270 0 0 CONDIODE
flabel metal1 s 362 3284 408 3414 0 FreeSans 200 0 0 0 PD_H
port 2 nsew
flabel metal1 s -50 2854 -7 2984 0 FreeSans 200 0 0 0 PAD
port 3 nsew
flabel metal1 s -50 4748 -7 4878 0 FreeSans 200 0 0 0 PAD
port 3 nsew
flabel metal1 s 362 4318 408 4448 0 FreeSans 200 0 0 0 PD_H
port 2 nsew
<< properties >>
string GDS_END 43339672
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43305116
<< end >>
