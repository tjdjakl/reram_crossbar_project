magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect -38 261 314 582
<< pwell >>
rect 1 21 275 177
rect 213 -17 247 21
<< scnmos >>
rect 79 47 109 151
rect 167 47 197 151
<< scpmoshvt >>
rect 79 339 109 497
rect 167 339 197 497
<< ndiff >>
rect 27 123 79 151
rect 27 89 35 123
rect 69 89 79 123
rect 27 47 79 89
rect 109 93 167 151
rect 109 59 121 93
rect 155 59 167 93
rect 109 47 167 59
rect 197 106 249 151
rect 197 72 207 106
rect 241 72 249 106
rect 197 47 249 72
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 396 79 443
rect 27 362 35 396
rect 69 362 79 396
rect 27 339 79 362
rect 109 477 167 497
rect 109 443 121 477
rect 155 443 167 477
rect 109 409 167 443
rect 109 375 121 409
rect 155 375 167 409
rect 109 339 167 375
rect 197 477 249 497
rect 197 443 207 477
rect 241 443 249 477
rect 197 409 249 443
rect 197 375 207 409
rect 241 375 249 409
rect 197 339 249 375
<< ndiffc >>
rect 35 89 69 123
rect 121 59 155 93
rect 207 72 241 106
<< pdiffc >>
rect 35 443 69 477
rect 35 362 69 396
rect 121 443 155 477
rect 121 375 155 409
rect 207 443 241 477
rect 207 375 241 409
<< poly >>
rect 79 497 109 523
rect 167 497 197 523
rect 79 278 109 339
rect 167 324 197 339
rect 167 300 203 324
rect 75 262 129 278
rect 75 228 85 262
rect 119 228 129 262
rect 75 212 129 228
rect 173 265 203 300
rect 173 249 249 265
rect 173 215 205 249
rect 239 215 249 249
rect 79 151 109 212
rect 173 199 249 215
rect 173 190 203 199
rect 167 166 203 190
rect 167 151 197 166
rect 79 21 109 47
rect 167 21 197 47
<< polycont >>
rect 85 228 119 262
rect 205 215 239 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 17 477 71 493
rect 17 443 35 477
rect 69 443 71 477
rect 17 396 71 443
rect 17 362 35 396
rect 69 362 71 396
rect 105 477 171 527
rect 105 443 121 477
rect 155 443 171 477
rect 105 409 171 443
rect 105 375 121 409
rect 155 375 171 409
rect 207 477 241 493
rect 207 409 241 443
rect 17 312 71 362
rect 207 341 241 375
rect 17 152 51 312
rect 108 307 241 341
rect 108 278 142 307
rect 85 262 142 278
rect 119 228 142 262
rect 85 212 142 228
rect 108 161 142 212
rect 189 249 255 271
rect 189 215 205 249
rect 239 215 255 249
rect 189 197 255 215
rect 17 123 69 152
rect 108 127 241 161
rect 17 89 35 123
rect 207 106 241 127
rect 17 51 69 89
rect 105 59 121 93
rect 155 59 171 93
rect 105 17 171 59
rect 207 51 241 72
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
flabel metal1 s 213 -17 247 17 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 213 527 247 561 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel locali s 29 85 63 119 0 FreeSans 200 180 0 0 X
port 6 nsew signal output
flabel locali s 29 357 63 391 0 FreeSans 200 180 0 0 X
port 6 nsew signal output
flabel locali s 29 425 63 459 0 FreeSans 200 180 0 0 X
port 6 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel nwell s 213 527 247 561 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 213 -17 247 17 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 clkbuf_1
rlabel metal1 s 0 -48 276 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 276 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 276 544
string GDS_END 3203066
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3199316
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 6.900 13.600 0.000 13.600 
<< end >>
