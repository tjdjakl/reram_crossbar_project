magic
tech sky130B
magscale 1 2
timestamp 1688980957
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 107 157 524 203
rect 1 21 827 157
rect 30 -17 64 21
<< locali >>
rect 17 212 111 325
rect 614 297 710 493
rect 671 128 710 297
rect 610 51 710 128
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 393 86 493
rect 120 427 186 527
rect 17 359 212 393
rect 178 249 212 359
rect 246 357 332 493
rect 366 393 420 493
rect 510 427 576 527
rect 366 358 580 393
rect 298 297 332 357
rect 178 215 264 249
rect 298 215 483 297
rect 546 249 580 358
rect 744 297 811 527
rect 546 215 637 249
rect 178 178 212 215
rect 298 181 332 215
rect 546 181 580 215
rect 17 144 212 178
rect 17 51 83 144
rect 117 17 183 110
rect 256 51 332 181
rect 366 147 580 181
rect 366 51 420 147
rect 510 17 576 113
rect 744 17 811 129
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 17 212 111 325 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 827 157 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 107 157 524 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 610 51 710 128 6 X
port 6 nsew signal output
rlabel locali s 671 128 710 297 6 X
port 6 nsew signal output
rlabel locali s 614 297 710 493 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3265580
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3259014
<< end >>
