magic
tech sky130B
magscale 1 2
timestamp 1700618825
<< pwell >>
rect -278 -333 278 333
<< mvnmos >>
rect -50 -75 50 75
<< mvndiff >>
rect -108 63 -50 75
rect -108 -63 -96 63
rect -62 -63 -50 63
rect -108 -75 -50 -63
rect 50 63 108 75
rect 50 -63 62 63
rect 96 -63 108 63
rect 50 -75 108 -63
<< mvndiffc >>
rect -96 -63 -62 63
rect 62 -63 96 63
<< mvpsubdiff >>
rect -242 285 242 297
rect -242 251 -134 285
rect 134 251 242 285
rect -242 239 242 251
rect -242 189 -184 239
rect -242 -189 -230 189
rect -196 -189 -184 189
rect 184 189 242 239
rect -242 -239 -184 -189
rect 184 -189 196 189
rect 230 -189 242 189
rect 184 -239 242 -189
rect -242 -251 242 -239
rect -242 -285 -134 -251
rect 134 -285 242 -251
rect -242 -297 242 -285
<< mvpsubdiffcont >>
rect -134 251 134 285
rect -230 -189 -196 189
rect 196 -189 230 189
rect -134 -285 134 -251
<< poly >>
rect -50 147 50 163
rect -50 113 -34 147
rect 34 113 50 147
rect -50 75 50 113
rect -50 -113 50 -75
rect -50 -147 -34 -113
rect 34 -147 50 -113
rect -50 -163 50 -147
<< polycont >>
rect -34 113 34 147
rect -34 -147 34 -113
<< locali >>
rect -230 251 -134 285
rect 134 251 230 285
rect -230 189 -196 251
rect 196 189 230 251
rect -50 113 -34 147
rect 34 113 50 147
rect -96 63 -62 79
rect -96 -79 -62 -63
rect 62 63 96 79
rect 62 -79 96 -63
rect -50 -147 -34 -113
rect 34 -147 50 -113
rect -230 -251 -196 -189
rect 196 -251 230 -189
rect -230 -285 -134 -251
rect 134 -285 230 -251
<< viali >>
rect -34 113 34 147
rect -96 -63 -62 63
rect 62 -63 96 63
rect -34 -147 34 -113
<< metal1 >>
rect -46 147 46 153
rect -46 113 -34 147
rect 34 113 46 147
rect -46 107 46 113
rect -102 63 -56 75
rect -102 -63 -96 63
rect -62 -63 -56 63
rect -102 -75 -56 -63
rect 56 63 102 75
rect 56 -63 62 63
rect 96 -63 102 63
rect 56 -75 102 -63
rect -46 -113 46 -107
rect -46 -147 -34 -113
rect 34 -147 46 -113
rect -46 -153 46 -147
<< properties >>
string FIXED_BBOX -213 -268 213 268
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.75 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
